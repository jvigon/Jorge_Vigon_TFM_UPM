use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_6_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_6_LAYER;

architecture Behavioral of ROM_FC_84_6_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_6: ROM_ARRAY_PESOS_FC_84 := (
"01011000", 
"01101110", 
"01110100", 
"10001111", 
"01111001", 
"01111001", 
"10100111", 
"10011000", 
"01101010", 
"01111101", 
"01110011", 
"00110011", 
"01110010", 
"01111010", 
"01100110", 
"10111111", 
"01101001", 
"10010011", 
"00111110", 
"10000110", 
"10011000", 
"01111100", 
"10101000", 
"01101110", 
"10001011", 
"01111101", 
"01011111", 
"10000100", 
"01010000", 
"01100100", 
"10001101", 
"01111001", 
"10010001", 
"01110110", 
"10010011", 
"10010100", 
"10110000", 
"01010010", 
"10011110", 
"10000111", 
"01101000", 
"01011100", 
"10011010", 
"10010011", 
"01011000", 
"01110110", 
"01010011", 
"01100111", 
"10000010", 
"10001110", 
"10000010", 
"01111001", 
"01110011", 
"01011011", 
"10000010", 
"01001111", 
"01110100", 
"01111001", 
"01110110", 
"01111001", 
"01011101", 
"10011111", 
"01101000", 
"01101001", 
"01011101", 
"01101111", 
"10110011", 
"10011000", 
"01100111", 
"01110001", 
"10000000", 
"01010010", 
"01100100", 
"01101100", 
"10001110", 
"10001100", 
"10010111", 
"10000111", 
"01110001", 
"01011010", 
"01101101", 
"01101011", 
"01101010", 
"01100110", 
"10001110", 
"01101110", 
"01101001", 
"01100111", 
"10000000", 
"10010111", 
"01100110", 
"10001001", 
"01010111", 
"01111011", 
"10011010", 
"01110001", 
"01111011", 
"10000000", 
"01111000", 
"10000000", 
"10000001", 
"01101110", 
"01111101", 
"00101100", 
"10000011", 
"01100101", 
"01111101", 
"01110010", 
"01101010", 
"10000001", 
"10000110", 
"10001001", 
"10001011", 
"10100111", 
"01110011", 
"01100001", 
"01111100", 
"01000110", 
"10000100", 
"01011111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_6 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_6(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
