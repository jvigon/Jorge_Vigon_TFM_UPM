use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_25_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_25_LAYER;

architecture Behavioral of ROM_FC_84_25_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_25: ROM_ARRAY_PESOS_FC_84 := (
"10000101", 
"10001011", 
"10010000", 
"01100111", 
"10010100", 
"10001100", 
"01111111", 
"01001110", 
"01111110", 
"01100100", 
"10101010", 
"10001001", 
"01111001", 
"01111000", 
"01111000", 
"01011100", 
"01111101", 
"10000001", 
"01101000", 
"01110011", 
"01011001", 
"01110000", 
"10000100", 
"01011010", 
"01111100", 
"10111001", 
"01101110", 
"01100011", 
"01001110", 
"01101100", 
"01110011", 
"01011110", 
"00111010", 
"10010111", 
"01110011", 
"10001011", 
"01100011", 
"01111101", 
"01110100", 
"01101011", 
"10010000", 
"10100001", 
"10001001", 
"01001101", 
"01100110", 
"01010110", 
"10001110", 
"01100010", 
"10001101", 
"01111110", 
"01100010", 
"01100111", 
"10000101", 
"10000001", 
"01011110", 
"01111000", 
"01101001", 
"10011000", 
"01101100", 
"10110010", 
"01110111", 
"01011000", 
"01100000", 
"01011001", 
"01101101", 
"10000000", 
"10000100", 
"01110100", 
"10011101", 
"01101010", 
"01111101", 
"10001000", 
"01101001", 
"10011001", 
"10001011", 
"01110000", 
"01111110", 
"10001100", 
"01101100", 
"10011110", 
"01100110", 
"01101001", 
"01110110", 
"01101100", 
"10000011", 
"01101010", 
"01100010", 
"01100110", 
"10011000", 
"10100000", 
"01011100", 
"10001011", 
"01011001", 
"01100111", 
"01111010", 
"10011000", 
"10001110", 
"10000110", 
"01011110", 
"01100000", 
"01100111", 
"10001011", 
"01010110", 
"00110101", 
"10100010", 
"10000000", 
"01111101", 
"01110111", 
"01010001", 
"10011100", 
"01110000", 
"10001001", 
"10001001", 
"10011111", 
"01110001", 
"10011101", 
"01011100", 
"10100001", 
"10001100", 
"10001011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_25 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_25(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
