use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_83_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_83_LAYER;

architecture Behavioral of ROM_FC_120_83_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_83: ROM_ARRAY_PESOS_FC_120 := (
"10000110", 
"10001110", 
"01110100", 
"10100011", 
"01110011", 
"10001010", 
"01101000", 
"10000101", 
"10000100", 
"00110101", 
"01000100", 
"10011011", 
"01100100", 
"10000111", 
"10000101", 
"10010001", 
"10010111", 
"10001100", 
"01101010", 
"01110000", 
"10001100", 
"10010010", 
"10001011", 
"10000011", 
"01110101", 
"01101111", 
"00110111", 
"01101100", 
"01101011", 
"01011101", 
"01111001", 
"01101010", 
"01111100", 
"01011101", 
"01001001", 
"01011011", 
"10010000", 
"11000010", 
"10100111", 
"01110001", 
"01110010", 
"01010110", 
"10001111", 
"10001100", 
"01001100", 
"01101100", 
"10010011", 
"10000000", 
"10001110", 
"01101010", 
"01111011", 
"10001110", 
"01111001", 
"10011110", 
"10110101", 
"01111000", 
"10000011", 
"10001011", 
"10000100", 
"10001010", 
"01000100", 
"10001110", 
"10000111", 
"10001110", 
"01111001", 
"10100100", 
"01001100", 
"01111100", 
"10011111", 
"10000111", 
"10001010", 
"10100100", 
"01110010", 
"10100111", 
"10100101", 
"10000100", 
"01110111", 
"01111011", 
"10000000", 
"01110110", 
"01110100", 
"10100011", 
"01010111", 
"01000000", 
"01100111", 
"01101101", 
"01011110", 
"01111111", 
"10011101", 
"01101110", 
"01000101", 
"10000101", 
"01101110", 
"01101001", 
"01111001", 
"10001100", 
"01111101", 
"01110100", 
"01001101", 
"01001111", 
"01110001", 
"10001111", 
"01110010", 
"10010110", 
"10001000", 
"01101100", 
"10011011", 
"10000101", 
"01011100", 
"01111000", 
"10000000", 
"01110111", 
"01111110", 
"00101111", 
"01111001", 
"10110001", 
"10000111", 
"01011010", 
"10011100", 
"10000100", 
"10011000", 
"10001110", 
"01110100", 
"01011011", 
"01001110", 
"10010111", 
"10010011", 
"01110011", 
"10010101", 
"01111010", 
"01011001", 
"10100001", 
"01111010", 
"01101011", 
"01101011", 
"10001110", 
"01111010", 
"10001011", 
"01110101", 
"01111010", 
"01001111", 
"01010101", 
"01111011", 
"01110010", 
"10010110", 
"01100011", 
"10101000", 
"10010000", 
"10000110", 
"10011000", 
"10000100", 
"01111011", 
"10100000", 
"01101101", 
"01011111", 
"01101011", 
"01001100", 
"01111010", 
"01110111", 
"01110100", 
"10110100", 
"00110000", 
"01110000", 
"10011000", 
"01110011", 
"10100100", 
"01001100", 
"01101001", 
"10001001", 
"01111010", 
"10001111", 
"10001111", 
"10001011", 
"10001111", 
"10001000", 
"01111100", 
"01110010", 
"00111100", 
"10100101", 
"11001111", 
"01110010", 
"10000001", 
"10010010", 
"01111000", 
"01111100", 
"10010010", 
"01111011", 
"10010000", 
"01001110", 
"01100001", 
"10000011", 
"10001100", 
"01111111", 
"10000001", 
"10011101", 
"01111111", 
"01111001", 
"10011001", 
"01111100", 
"10000111", 
"10001101", 
"10011001", 
"01101110", 
"10001011", 
"10000110", 
"00101011", 
"01101111", 
"01111111", 
"10100000", 
"01100001", 
"10011101", 
"01100000", 
"10000010", 
"10100010", 
"00111000", 
"01010001", 
"01111101", 
"10001000", 
"10100011", 
"10011110", 
"10001010", 
"01101110", 
"01101110", 
"10000111", 
"10000101", 
"01001110", 
"10000100", 
"10001001", 
"10001110", 
"01111100", 
"01101101", 
"01101010", 
"01110100", 
"10010010", 
"10100101", 
"11000100", 
"01111011", 
"10011000", 
"10000100", 
"01111111", 
"00111010", 
"01011011", 
"01110111", 
"10011111", 
"10001010", 
"01011011", 
"10000010", 
"01010101", 
"10000011", 
"10000101", 
"10010011", 
"10010011", 
"01100111", 
"01110100", 
"10001110", 
"01111101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_83: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_83(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
