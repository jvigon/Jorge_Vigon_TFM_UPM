use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_10_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_10_LAYER;

architecture Behavioral of ROM_FC_84_10_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_10: ROM_ARRAY_PESOS_FC_84 := (
"01111000", 
"01001110", 
"00110101", 
"10010101", 
"10100001", 
"10001111", 
"10010111", 
"01101001", 
"10100011", 
"01111001", 
"10001001", 
"01111100", 
"01000100", 
"10010000", 
"01111110", 
"01111001", 
"01110110", 
"01101001", 
"01011111", 
"01111011", 
"10011011", 
"01000010", 
"10100000", 
"01011010", 
"01111111", 
"10111010", 
"01111001", 
"01100110", 
"01100001", 
"10000111", 
"10010010", 
"10001011", 
"01011011", 
"10001001", 
"01011101", 
"10001101", 
"01100110", 
"01010001", 
"10011111", 
"10100000", 
"01100110", 
"01111010", 
"10010110", 
"01110101", 
"01011110", 
"01111100", 
"10011001", 
"01010000", 
"01111001", 
"10011100", 
"01101011", 
"01101001", 
"01110010", 
"01111111", 
"01100111", 
"10100011", 
"01110100", 
"10010001", 
"01111111", 
"01100100", 
"01111100", 
"10010110", 
"10001001", 
"01000110", 
"10110100", 
"01101100", 
"01100000", 
"01111011", 
"10000100", 
"01001101", 
"01010100", 
"10001100", 
"10000000", 
"10010110", 
"10000010", 
"10001000", 
"10000111", 
"10001110", 
"01110101", 
"10000110", 
"10011000", 
"01111101", 
"01000000", 
"01010110", 
"10100000", 
"10000001", 
"01011010", 
"10010000", 
"01101001", 
"10011110", 
"00111101", 
"10000010", 
"01111010", 
"10001000", 
"01011000", 
"10001111", 
"10000011", 
"10100001", 
"01000100", 
"10001010", 
"01111010", 
"10000100", 
"01000000", 
"01100111", 
"01110001", 
"10001100", 
"01101110", 
"01100110", 
"10000000", 
"11000101", 
"01111010", 
"01101011", 
"10010010", 
"01101000", 
"01101101", 
"10011001", 
"10000001", 
"10111111", 
"01101101", 
"01011101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_10 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_10(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
