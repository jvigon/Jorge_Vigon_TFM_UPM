use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_16_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_16_LAYER;

architecture Behavioral of ROM_FC_120_16_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_16: ROM_ARRAY_PESOS_FC_120 := (
"01101111", 
"01110110", 
"10000000", 
"01001100", 
"10010010", 
"01000110", 
"01111101", 
"10010101", 
"10000001", 
"10100101", 
"10011111", 
"01110010", 
"10011101", 
"01010101", 
"01111010", 
"01101111", 
"01111110", 
"01110010", 
"10000110", 
"00111101", 
"10000001", 
"01011110", 
"01110100", 
"10010011", 
"01101011", 
"01111101", 
"10000110", 
"10100000", 
"10010011", 
"01010110", 
"10001100", 
"01111101", 
"01100001", 
"10001100", 
"01110110", 
"01110101", 
"01110001", 
"01101111", 
"01110000", 
"01011001", 
"01110010", 
"01110000", 
"01111100", 
"01111111", 
"10001101", 
"10010101", 
"01110110", 
"10011110", 
"10000111", 
"10010101", 
"01110011", 
"10101010", 
"10000000", 
"10010100", 
"10001001", 
"01011001", 
"01101101", 
"01000110", 
"10000000", 
"00111100", 
"10011110", 
"10001100", 
"10010011", 
"10010001", 
"10001100", 
"01110101", 
"01111001", 
"10100111", 
"10010111", 
"10010111", 
"01101010", 
"10011001", 
"01101001", 
"01011001", 
"01111010", 
"10000001", 
"01111001", 
"10010001", 
"01111000", 
"10000111", 
"01110110", 
"01110100", 
"01100111", 
"01110100", 
"01110111", 
"10000101", 
"01011001", 
"01101100", 
"01110111", 
"01101010", 
"10001000", 
"01101111", 
"01101101", 
"01111001", 
"01111111", 
"10010111", 
"01100010", 
"10101000", 
"10010110", 
"01111010", 
"10000011", 
"01100100", 
"01100010", 
"01101001", 
"01111010", 
"01110110", 
"10000100", 
"10000000", 
"01100011", 
"01100101", 
"01111111", 
"01111001", 
"01101101", 
"10000000", 
"10001101", 
"10011100", 
"10000000", 
"10010001", 
"01111110", 
"10011111", 
"01101011", 
"01011110", 
"01111111", 
"01110001", 
"01101101", 
"01100011", 
"10010101", 
"01011001", 
"10001101", 
"01100001", 
"01111010", 
"01110001", 
"01100100", 
"10011110", 
"00111111", 
"01110010", 
"01111001", 
"01010111", 
"01011111", 
"01100011", 
"01100001", 
"11010000", 
"01110010", 
"01111011", 
"01110010", 
"01010011", 
"01011001", 
"10000110", 
"01101100", 
"10001010", 
"01101111", 
"01110010", 
"01101011", 
"01111101", 
"01110001", 
"01100101", 
"01111110", 
"10100100", 
"10000011", 
"01100101", 
"01011100", 
"01101100", 
"10010110", 
"01111000", 
"01110000", 
"10010010", 
"10001111", 
"01110101", 
"01111111", 
"01001001", 
"01011111", 
"10001011", 
"10011110", 
"10000011", 
"10000111", 
"10000100", 
"01111000", 
"10011101", 
"01001111", 
"01011111", 
"10010100", 
"10010000", 
"10100110", 
"01101101", 
"01101111", 
"01011110", 
"01110010", 
"01010110", 
"01110101", 
"10100101", 
"10001110", 
"10000011", 
"01111011", 
"10001000", 
"10001110", 
"10011001", 
"10001001", 
"10101001", 
"01111101", 
"10001010", 
"10010001", 
"01100110", 
"10000011", 
"10000101", 
"10100001", 
"10011001", 
"01101111", 
"01101110", 
"01110101", 
"01010111", 
"01110101", 
"01010111", 
"01110110", 
"01110101", 
"11000100", 
"10100001", 
"01101110", 
"01110001", 
"01111110", 
"10001001", 
"10001001", 
"10000011", 
"01111111", 
"01110010", 
"10001100", 
"01111010", 
"01011110", 
"01100111", 
"01110100", 
"01101110", 
"01111010", 
"01110101", 
"01111000", 
"10001011", 
"01010011", 
"01111010", 
"10100110", 
"10011001", 
"10010011", 
"01110100", 
"10001011", 
"01111110", 
"01110011", 
"01101101", 
"10010110", 
"10100000", 
"10000000", 
"10011000", 
"10000101", 
"10011101", 
"01110010", 
"01010000", 
"01111000", 
"01001110", 
"01111101", 
"10000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_16: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_16(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
