use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_103_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_103_LAYER;

architecture Behavioral of ROM_FC_120_103_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_103: ROM_ARRAY_PESOS_FC_120 := (
"01110100", 
"10000010", 
"01111100", 
"01011111", 
"01101010", 
"01001111", 
"00000000", 
"00110100", 
"10000101", 
"10011000", 
"10111010", 
"10100100", 
"01111110", 
"11000101", 
"10001111", 
"01101101", 
"01000111", 
"10000111", 
"01100100", 
"01011000", 
"01101111", 
"01011010", 
"00111101", 
"01110111", 
"01110110", 
"10010000", 
"10000111", 
"10110001", 
"10010001", 
"01111110", 
"10101011", 
"10011010", 
"01011010", 
"10010001", 
"01010001", 
"01000101", 
"10001110", 
"10001100", 
"01101011", 
"01100001", 
"01111000", 
"01101100", 
"01101001", 
"10011111", 
"10001110", 
"01101000", 
"10000101", 
"01111100", 
"10100111", 
"11010100", 
"01101101", 
"10001111", 
"01101011", 
"10001011", 
"10001100", 
"01101101", 
"10000011", 
"01010010", 
"10100100", 
"10000110", 
"01110110", 
"01111011", 
"01111111", 
"10000011", 
"01111011", 
"01010110", 
"01101011", 
"00100101", 
"01011001", 
"01100110", 
"01001011", 
"10000111", 
"01110011", 
"01111010", 
"01011001", 
"10111101", 
"10001000", 
"10100001", 
"10000010", 
"10001111", 
"01110001", 
"01111111", 
"10001010", 
"00001001", 
"01101000", 
"01110010", 
"01101010", 
"01110111", 
"10001111", 
"01111011", 
"01110101", 
"10101101", 
"11000010", 
"01100110", 
"10011101", 
"10000111", 
"01110100", 
"01011101", 
"10001001", 
"01011101", 
"01010111", 
"10000111", 
"01100011", 
"10110100", 
"10010010", 
"10001110", 
"01110100", 
"10100001", 
"10101001", 
"00111010", 
"10001100", 
"10010110", 
"01101000", 
"01110110", 
"10000100", 
"10110101", 
"01110001", 
"01111111", 
"01010100", 
"10101111", 
"01010101", 
"01111111", 
"10100110", 
"01111101", 
"10000001", 
"01011101", 
"01111111", 
"10000101", 
"01101011", 
"01010011", 
"10010101", 
"10001000", 
"00010110", 
"01100100", 
"01101010", 
"01000001", 
"01101011", 
"01001011", 
"01001101", 
"01100011", 
"01111101", 
"10110010", 
"10010000", 
"10001000", 
"01010001", 
"01010111", 
"10001010", 
"01101011", 
"10100001", 
"01100001", 
"01101100", 
"01111001", 
"01101110", 
"10100100", 
"01100101", 
"01111100", 
"10101000", 
"10101010", 
"10100100", 
"01111011", 
"01000111", 
"01111001", 
"10011000", 
"10000100", 
"01111010", 
"01111001", 
"01000111", 
"01101001", 
"01110001", 
"01111001", 
"10100100", 
"01011010", 
"01100000", 
"00111111", 
"10001100", 
"10011000", 
"01100101", 
"10100011", 
"01111000", 
"01101100", 
"01111000", 
"01101111", 
"01111101", 
"01100110", 
"10000111", 
"10000111", 
"10001001", 
"01101110", 
"10011000", 
"10010001", 
"10111110", 
"10010110", 
"01100001", 
"10100011", 
"10101110", 
"01101100", 
"00110110", 
"10101000", 
"10100100", 
"01100111", 
"10001000", 
"01111110", 
"10101010", 
"10001010", 
"10011011", 
"11011110", 
"10100111", 
"01111011", 
"10001011", 
"10010011", 
"01101001", 
"01111110", 
"01111111", 
"01110001", 
"10100000", 
"01100011", 
"10101011", 
"01110101", 
"10011000", 
"10000010", 
"10100011", 
"10101111", 
"11000100", 
"10011111", 
"10010101", 
"10010000", 
"01010000", 
"10001001", 
"10100111", 
"10000100", 
"10011011", 
"10010001", 
"10010010", 
"10000011", 
"10010001", 
"01000110", 
"01101010", 
"10000011", 
"01111011", 
"01111010", 
"01111010", 
"10100000", 
"00111001", 
"01011111", 
"10001011", 
"10011111", 
"10001110", 
"10101110", 
"01111001", 
"01101001", 
"10100110", 
"01100110", 
"01010101", 
"01111110", 
"01100000", 
"01110011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_103 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_103(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
