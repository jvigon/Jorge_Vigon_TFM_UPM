use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_23_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_23_LAYER;

architecture Behavioral of ROM_FC_120_23_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_23: ROM_ARRAY_PESOS_FC_120 := (
"10000010", 
"01101011", 
"10001100", 
"01101100", 
"01010111", 
"01100010", 
"10000110", 
"01000110", 
"01100111", 
"10011000", 
"10101101", 
"01001100", 
"10011111", 
"01100101", 
"10001011", 
"10010001", 
"10011011", 
"10000101", 
"01100111", 
"01010010", 
"10000010", 
"10000111", 
"01001111", 
"10000010", 
"01101000", 
"10001001", 
"10001001", 
"01110000", 
"10001010", 
"10001111", 
"10011001", 
"10001111", 
"01010111", 
"01110101", 
"01110011", 
"01111001", 
"10000100", 
"10011000", 
"01010111", 
"10010111", 
"01110100", 
"01101001", 
"01110010", 
"01100100", 
"01110110", 
"10110110", 
"10001001", 
"10000100", 
"01111111", 
"01110010", 
"01011000", 
"01111100", 
"01110011", 
"10011110", 
"10000110", 
"01000110", 
"01110001", 
"01101101", 
"01101000", 
"01110110", 
"10010100", 
"10011110", 
"10001100", 
"01111111", 
"10011001", 
"10001111", 
"01010000", 
"01010101", 
"01110101", 
"10010010", 
"01100010", 
"01101111", 
"01110001", 
"10000110", 
"10100011", 
"10001101", 
"01101010", 
"00011110", 
"01111010", 
"01100110", 
"01101100", 
"10101110", 
"01100001", 
"01011000", 
"01110111", 
"01011011", 
"10011101", 
"10001011", 
"01101101", 
"01011100", 
"10010111", 
"01110001", 
"10000101", 
"10010000", 
"10000010", 
"01110010", 
"10001110", 
"01110111", 
"01110100", 
"01111100", 
"10000011", 
"01111000", 
"01111000", 
"01010001", 
"01111110", 
"10000001", 
"01011100", 
"01110001", 
"01011011", 
"10010010", 
"10000000", 
"10010011", 
"10100001", 
"10001011", 
"01101001", 
"01111110", 
"10001100", 
"01101101", 
"00111000", 
"10100110", 
"10010011", 
"10110011", 
"10001100", 
"01110011", 
"01011100", 
"01101001", 
"10000101", 
"10001011", 
"10010001", 
"01100001", 
"00101101", 
"01010000", 
"10101000", 
"10000001", 
"10110100", 
"10111111", 
"10001000", 
"01011000", 
"01000011", 
"10111001", 
"10010111", 
"01101011", 
"10010000", 
"10000010", 
"01111111", 
"10011000", 
"01110101", 
"01011010", 
"10001111", 
"01011111", 
"10110000", 
"01101101", 
"01111010", 
"00101001", 
"00111011", 
"01100110", 
"10110110", 
"10100011", 
"01110010", 
"10000000", 
"10010110", 
"01100011", 
"01101010", 
"01011111", 
"10001101", 
"10000000", 
"01100111", 
"10000100", 
"10000011", 
"01010010", 
"10011000", 
"01101110", 
"10000111", 
"01110011", 
"10010010", 
"01111010", 
"01111100", 
"01100111", 
"01110010", 
"10011100", 
"01111011", 
"10000001", 
"01100111", 
"10100101", 
"10000001", 
"01100001", 
"10000010", 
"01011100", 
"00110111", 
"01110111", 
"01110000", 
"01110101", 
"01100011", 
"01100010", 
"10011111", 
"01101000", 
"10011001", 
"10001111", 
"10010011", 
"01011001", 
"01110111", 
"01011111", 
"01101101", 
"10001010", 
"10000101", 
"01011101", 
"10000100", 
"01111100", 
"01100110", 
"10100000", 
"01111001", 
"01111101", 
"10010000", 
"01111100", 
"10000100", 
"01001010", 
"01011111", 
"01010100", 
"10000110", 
"01011001", 
"01110011", 
"01001010", 
"01110000", 
"10000000", 
"10000100", 
"01110111", 
"01110000", 
"10001010", 
"10001111", 
"10100101", 
"01100011", 
"01110111", 
"10100001", 
"01100101", 
"11000001", 
"01100111", 
"10010111", 
"01110011", 
"10001001", 
"10000011", 
"01110000", 
"10010111", 
"00101011", 
"01010010", 
"10001111", 
"10011110", 
"10100110", 
"01110011", 
"01110100", 
"01001100", 
"10000101", 
"01010110", 
"01110111", 
"10101001", 
"01110011", 
"01111000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_23: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_23(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
