use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_22_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_22_LAYER;

architecture Behavioral of ROM_FC_84_22_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_22: ROM_ARRAY_PESOS_FC_84 := (
"10000100", 
"10001010", 
"01100101", 
"01110110", 
"01111011", 
"10010010", 
"10000000", 
"01010111", 
"10000101", 
"01111100", 
"10001011", 
"01101000", 
"10001000", 
"10001010", 
"01000111", 
"01101011", 
"01110100", 
"10001100", 
"01101001", 
"01111111", 
"01001110", 
"01010011", 
"01111011", 
"10101100", 
"10000110", 
"10001101", 
"10101000", 
"10010001", 
"10011100", 
"01010100", 
"01110011", 
"00111111", 
"10001000", 
"10000010", 
"10011000", 
"01100010", 
"10100011", 
"10110000", 
"01011000", 
"01011111", 
"01101110", 
"01001101", 
"10000101", 
"10001111", 
"01011010", 
"01110100", 
"10100010", 
"01110001", 
"01111001", 
"10001100", 
"01111111", 
"10001100", 
"01110101", 
"10001111", 
"01101000", 
"10001111", 
"10000100", 
"01110010", 
"01101101", 
"10010111", 
"01101111", 
"01000110", 
"10101001", 
"10111000", 
"01111100", 
"01110111", 
"10011100", 
"10011110", 
"01110110", 
"01101011", 
"10101101", 
"00110011", 
"10011111", 
"10010010", 
"10100111", 
"01111100", 
"10000110", 
"10000010", 
"10000011", 
"01100011", 
"10001000", 
"01100100", 
"10011000", 
"01101110", 
"01010110", 
"10010010", 
"01110001", 
"10100100", 
"01110011", 
"01110001", 
"10010000", 
"10100100", 
"01100101", 
"01001111", 
"10001010", 
"10011000", 
"10010111", 
"10001100", 
"01100101", 
"01111010", 
"01110011", 
"10010110", 
"01101010", 
"10000110", 
"10000011", 
"10000100", 
"01110000", 
"10010101", 
"01100000", 
"10011010", 
"00110000", 
"10000111", 
"10001000", 
"01101100", 
"10010101", 
"10011001", 
"01101101", 
"10010010", 
"01100110", 
"10101111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_22 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_22(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
