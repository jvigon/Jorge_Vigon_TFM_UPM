use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_9_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_9_LAYER;

architecture Behavioral of ROM_FC_120_9_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_9: ROM_ARRAY_PESOS_FC_120 := (
"01011001", 
"01100000", 
"10000100", 
"10001010", 
"01001100", 
"01100001", 
"01011001", 
"01101001", 
"01111000", 
"10001010", 
"01110011", 
"01001010", 
"01100101", 
"00101010", 
"10001101", 
"10000011", 
"01110101", 
"01110000", 
"10000110", 
"01110111", 
"10110101", 
"01000100", 
"01111111", 
"01100011", 
"10001001", 
"01100000", 
"01111001", 
"10011101", 
"01101011", 
"01111011", 
"10000000", 
"01111111", 
"01011011", 
"01011100", 
"01101110", 
"01111011", 
"10010001", 
"01010000", 
"01000100", 
"01110000", 
"01110100", 
"10110001", 
"01101001", 
"10011100", 
"10000000", 
"01010010", 
"01111111", 
"10001001", 
"01110001", 
"01100101", 
"01100111", 
"01100000", 
"01100000", 
"10000000", 
"01111000", 
"01010101", 
"01101110", 
"10001011", 
"01101011", 
"01111100", 
"01011011", 
"00111011", 
"10001010", 
"10001000", 
"01101001", 
"01111000", 
"01011000", 
"10000011", 
"01010111", 
"01100111", 
"01100010", 
"01111011", 
"01110100", 
"01110000", 
"01011100", 
"01011111", 
"01001010", 
"10110000", 
"01110000", 
"10010010", 
"01011101", 
"01110001", 
"01100010", 
"01101100", 
"01110110", 
"01100100", 
"10001100", 
"01110001", 
"01110000", 
"01011101", 
"01111011", 
"01110001", 
"01011110", 
"10001100", 
"01111101", 
"10000101", 
"01100011", 
"01101010", 
"01100010", 
"10100011", 
"01111110", 
"01101010", 
"01110110", 
"10001000", 
"10000001", 
"01100101", 
"01111011", 
"01101100", 
"10000001", 
"01011000", 
"01101101", 
"10001010", 
"01111000", 
"00110010", 
"10001100", 
"01111001", 
"10000000", 
"01100101", 
"01011110", 
"01100011", 
"01101101", 
"10001000", 
"01101101", 
"01111100", 
"01010101", 
"10001000", 
"10000111", 
"10000110", 
"01101100", 
"01101101", 
"01010010", 
"01011100", 
"10010000", 
"01110010", 
"10110011", 
"10110111", 
"10001010", 
"01101110", 
"01010111", 
"10010011", 
"01111011", 
"00010011", 
"10010000", 
"10010000", 
"10000000", 
"10000011", 
"01100010", 
"01011010", 
"10100001", 
"01001011", 
"10010110", 
"01011100", 
"10001111", 
"01001011", 
"01000001", 
"01011001", 
"10000011", 
"01100001", 
"10000111", 
"10000100", 
"10010101", 
"10000010", 
"01110111", 
"01011010", 
"01111111", 
"01010101", 
"01111110", 
"01001010", 
"10010010", 
"01011111", 
"10011100", 
"01100000", 
"01101111", 
"10001101", 
"10001001", 
"01111101", 
"01100101", 
"10010000", 
"01100110", 
"01100011", 
"01110100", 
"01110011", 
"01101010", 
"00111000", 
"01111111", 
"01011011", 
"01110000", 
"01110100", 
"01100110", 
"00110100", 
"10000111", 
"01110010", 
"01110010", 
"01101111", 
"10010110", 
"01101110", 
"10100101", 
"01100010", 
"01011010", 
"10000010", 
"01110111", 
"01111111", 
"01111001", 
"01111111", 
"10001010", 
"01101011", 
"01111011", 
"01101010", 
"01110110", 
"10000100", 
"10001011", 
"01100001", 
"01010011", 
"10001101", 
"01110011", 
"10010011", 
"01111101", 
"10001110", 
"01101100", 
"10000010", 
"10001101", 
"01100101", 
"01110011", 
"10010100", 
"10000110", 
"01111110", 
"01011111", 
"01000111", 
"01110001", 
"01011110", 
"01110101", 
"10101011", 
"01110100", 
"01100000", 
"01100001", 
"10001101", 
"01111011", 
"00111110", 
"01110011", 
"01101100", 
"01111101", 
"01100101", 
"10000101", 
"01110100", 
"01111100", 
"01010010", 
"10000000", 
"10000100", 
"01101110", 
"01110000", 
"01001011", 
"01101110", 
"01010111", 
"10011010", 
"10000101", 
"10010101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_9 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_9(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
