use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_54_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_54_LAYER;

architecture Behavioral of ROM_FC_120_54_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_54: ROM_ARRAY_PESOS_FC_120 := (
"10100000", 
"01100011", 
"01010011", 
"10010001", 
"01100011", 
"01101011", 
"01000010", 
"01100011", 
"01111111", 
"01010101", 
"01101101", 
"01001101", 
"01010010", 
"01100111", 
"10000111", 
"01101101", 
"10010001", 
"10010010", 
"01100100", 
"01101001", 
"01001010", 
"01111000", 
"10010001", 
"10101010", 
"01111010", 
"01101011", 
"01001000", 
"00100101", 
"01000101", 
"01101001", 
"01101011", 
"01101010", 
"10001011", 
"00110101", 
"01101101", 
"00110111", 
"01111011", 
"10110001", 
"10011011", 
"10100101", 
"01101111", 
"10000001", 
"10001110", 
"01110111", 
"01110111", 
"10011001", 
"10000110", 
"10010100", 
"10001000", 
"01110101", 
"10011100", 
"10010101", 
"10001001", 
"10011011", 
"01101010", 
"10010101", 
"01110000", 
"01111010", 
"10010011", 
"10010011", 
"10001000", 
"10100001", 
"01110000", 
"10000111", 
"10001011", 
"10010000", 
"01101111", 
"10010110", 
"01010111", 
"01101101", 
"01100101", 
"10101010", 
"01111001", 
"01100111", 
"10000010", 
"01100110", 
"01111101", 
"10101100", 
"10010000", 
"10001101", 
"01011100", 
"10000110", 
"01100100", 
"01101111", 
"01001100", 
"01101011", 
"10000000", 
"10000110", 
"10001101", 
"01001100", 
"01001001", 
"01100001", 
"10011100", 
"01100100", 
"10001011", 
"10001101", 
"10101001", 
"01110010", 
"01011011", 
"00011010", 
"10000110", 
"01111011", 
"10001011", 
"01111111", 
"10010010", 
"10011101", 
"10001110", 
"01011110", 
"01101101", 
"01001100", 
"01111100", 
"01111001", 
"01111100", 
"00111010", 
"10000001", 
"01111110", 
"10010010", 
"01011110", 
"01111101", 
"10000101", 
"01110100", 
"10101111", 
"10011010", 
"10010000", 
"10000100", 
"01111000", 
"10001011", 
"10001001", 
"01110011", 
"01111101", 
"01100110", 
"01111100", 
"01101010", 
"10000001", 
"01110001", 
"10011011", 
"10010000", 
"10010100", 
"01111100", 
"01110111", 
"01110100", 
"01011101", 
"10000110", 
"01101111", 
"10100101", 
"10001000", 
"01101101", 
"01111100", 
"01111110", 
"10111001", 
"10000001", 
"10000001", 
"01111010", 
"10010001", 
"01011111", 
"01110000", 
"10000000", 
"01110011", 
"01111001", 
"01111110", 
"10110101", 
"10010100", 
"01100110", 
"01100000", 
"10000101", 
"10011011", 
"10001010", 
"01111100", 
"01111011", 
"01111011", 
"10100011", 
"01100001", 
"01011100", 
"10101011", 
"01110011", 
"10001101", 
"01100001", 
"01110111", 
"10011011", 
"01010101", 
"01110010", 
"01100011", 
"01100001", 
"01111001", 
"10001001", 
"01101000", 
"01100101", 
"10100000", 
"01101100", 
"01011110", 
"10000001", 
"10000101", 
"01110100", 
"10101001", 
"10010001", 
"01010111", 
"01110101", 
"10111111", 
"01011100", 
"01101110", 
"01110100", 
"10000000", 
"01110101", 
"10100010", 
"10001101", 
"01100010", 
"10001000", 
"01101111", 
"10011111", 
"10001110", 
"01010011", 
"01001101", 
"01110001", 
"10111000", 
"01101010", 
"10110100", 
"01111000", 
"10000011", 
"10011001", 
"01110111", 
"10100100", 
"01001011", 
"01110010", 
"01111110", 
"01010111", 
"01000011", 
"01101101", 
"10010011", 
"01111010", 
"01111000", 
"01100001", 
"10010110", 
"01011111", 
"01110001", 
"10001101", 
"10000110", 
"01111100", 
"11010111", 
"10000111", 
"01110100", 
"01000011", 
"01111100", 
"10000100", 
"00111000", 
"10000000", 
"01100000", 
"10100100", 
"01101101", 
"10000111", 
"01101001", 
"01100111", 
"01100111", 
"01100001", 
"01101001", 
"10000111", 
"01110001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_54: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_54(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
