use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_98_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_98_LAYER;

architecture Behavioral of ROM_FC_120_98_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_98: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"01100110", 
"00110000", 
"01010110", 
"10011111", 
"01110010", 
"10101001", 
"10000111", 
"01110011", 
"10001111", 
"01111111", 
"10010011", 
"10010001", 
"01100010", 
"01111010", 
"10001010", 
"10010011", 
"01110011", 
"01101010", 
"00111101", 
"10000010", 
"10011110", 
"01101101", 
"01101000", 
"01110010", 
"01111101", 
"10001001", 
"01101000", 
"10110101", 
"01010011", 
"01111011", 
"01111010", 
"01111000", 
"01011110", 
"01001110", 
"01101110", 
"01101000", 
"01100010", 
"01011100", 
"01110001", 
"01110001", 
"10100000", 
"01110111", 
"10001101", 
"10011011", 
"10000010", 
"01111110", 
"01110011", 
"01110100", 
"01011011", 
"01101011", 
"01011000", 
"10001011", 
"01111100", 
"01100000", 
"01101100", 
"10001001", 
"10011010", 
"01011010", 
"01100111", 
"10000100", 
"01110101", 
"01110111", 
"01100110", 
"01110110", 
"01110111", 
"00111101", 
"00110110", 
"10001101", 
"10110000", 
"01101111", 
"01011100", 
"10001010", 
"01100100", 
"10101011", 
"01000111", 
"01100110", 
"10001010", 
"01111110", 
"01111000", 
"10001000", 
"10001010", 
"01101100", 
"10011011", 
"10001110", 
"01010100", 
"10000101", 
"10000101", 
"10001000", 
"01001110", 
"10001100", 
"00101100", 
"01100001", 
"10100010", 
"10000000", 
"10000011", 
"01110010", 
"01110001", 
"10100110", 
"10011011", 
"01110010", 
"01101111", 
"10011011", 
"10001101", 
"10010100", 
"10000010", 
"01101100", 
"01010111", 
"01100010", 
"01110101", 
"01110010", 
"01110100", 
"10010110", 
"01110000", 
"01110001", 
"01010101", 
"10001010", 
"10011110", 
"01010111", 
"01111010", 
"10001001", 
"10101010", 
"10001010", 
"10100101", 
"01111011", 
"01011110", 
"10000000", 
"10000100", 
"10001000", 
"10001111", 
"01110111", 
"11000010", 
"10100010", 
"01110111", 
"10001110", 
"01000100", 
"10001011", 
"00101011", 
"01011101", 
"10001111", 
"10000001", 
"11001110", 
"01111111", 
"10010100", 
"01100011", 
"01110001", 
"10000000", 
"11000000", 
"10001011", 
"01000100", 
"10010011", 
"01110111", 
"10010000", 
"01100011", 
"01110000", 
"01001001", 
"10000100", 
"10010111", 
"10001110", 
"10010001", 
"10000001", 
"01110101", 
"01010010", 
"01110000", 
"01110100", 
"10001001", 
"10010010", 
"01111000", 
"01111101", 
"10001000", 
"01111010", 
"01100100", 
"01110100", 
"10000101", 
"01101110", 
"10000101", 
"01111010", 
"01001110", 
"01110110", 
"10001001", 
"10001100", 
"10010001", 
"00100011", 
"10101000", 
"01110111", 
"10101010", 
"10001110", 
"10011000", 
"00000110", 
"01001000", 
"10000001", 
"10000111", 
"10000100", 
"10000001", 
"01011101", 
"01100111", 
"10100010", 
"01110010", 
"01110111", 
"01100111", 
"01101100", 
"01110110", 
"01011011", 
"10001001", 
"10101011", 
"01111011", 
"10000001", 
"10010000", 
"01011010", 
"10101100", 
"10001001", 
"01110111", 
"01110111", 
"10000110", 
"01010100", 
"01101010", 
"10001010", 
"01101010", 
"10111000", 
"10001010", 
"01110011", 
"01111101", 
"10010000", 
"10001001", 
"01101001", 
"10000110", 
"01000110", 
"01010001", 
"10001000", 
"10101010", 
"01111000", 
"01110000", 
"10000110", 
"01100100", 
"10011111", 
"01001110", 
"01101011", 
"01111010", 
"10000111", 
"10001100", 
"10000110", 
"01110110", 
"01101011", 
"00111010", 
"01110010", 
"10010100", 
"01110111", 
"01101000", 
"01110001", 
"01100100", 
"10100000", 
"01010010", 
"00111101", 
"10010100", 
"01111100", 
"10001101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_98: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_98(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
