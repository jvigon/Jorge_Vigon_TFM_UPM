use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_27_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_27_LAYER;

architecture Behavioral of ROM_FC_84_27_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_27: ROM_ARRAY_PESOS_FC_84 := (
"01001001", 
"10000110", 
"01110101", 
"10001011", 
"01110111", 
"01100100", 
"10010110", 
"01000000", 
"01001100", 
"01011111", 
"01101111", 
"01111100", 
"10100100", 
"01010010", 
"01010001", 
"10001100", 
"10001010", 
"01110011", 
"10010011", 
"10000101", 
"10010110", 
"10011110", 
"01101011", 
"10001010", 
"01111101", 
"01110101", 
"10000101", 
"01101000", 
"01101110", 
"01100011", 
"01110000", 
"00111011", 
"01010111", 
"01100010", 
"01001011", 
"01100010", 
"10011100", 
"10000111", 
"01101010", 
"10010010", 
"01110100", 
"01100110", 
"01111011", 
"10001010", 
"01110111", 
"01001100", 
"01011100", 
"10011101", 
"01101001", 
"01111001", 
"01110011", 
"01110010", 
"10001111", 
"01111110", 
"10001001", 
"10001001", 
"10010100", 
"01110111", 
"01111111", 
"10110101", 
"01100010", 
"10011011", 
"01110100", 
"01110000", 
"01011000", 
"01011001", 
"01100110", 
"10010100", 
"01111111", 
"01110100", 
"01100100", 
"01111001", 
"01111001", 
"01101000", 
"01111010", 
"01111000", 
"10101000", 
"10010111", 
"10000001", 
"10010111", 
"01010111", 
"01010110", 
"10001000", 
"01111000", 
"01011100", 
"01110100", 
"10100110", 
"10000110", 
"01111101", 
"10000100", 
"01110110", 
"01101000", 
"10101000", 
"10110100", 
"01101111", 
"01111010", 
"10001101", 
"10010000", 
"01101001", 
"10001011", 
"10010000", 
"10101100", 
"10000101", 
"10011001", 
"10010001", 
"10011000", 
"10000000", 
"01101010", 
"01010110", 
"01011000", 
"01010110", 
"01110111", 
"10011000", 
"10011101", 
"01101100", 
"01111011", 
"01100011", 
"10100111", 
"10011000", 
"01101010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_27 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_27(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
