use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_12_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_12_LAYER;

architecture Behavioral of ROM_FC_120_12_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_12: ROM_ARRAY_PESOS_FC_120 := (
"01111110", 
"10101111", 
"10010001", 
"10100010", 
"01101111", 
"10011011", 
"01110010", 
"10000100", 
"01111100", 
"10111010", 
"10011011", 
"01010101", 
"01111001", 
"10001111", 
"10001111", 
"10000010", 
"10001001", 
"10001100", 
"10000000", 
"01111111", 
"10000011", 
"10101110", 
"01111100", 
"01101011", 
"10000110", 
"10010001", 
"01101110", 
"10001011", 
"01011100", 
"11000101", 
"01110111", 
"10100011", 
"10001111", 
"10010110", 
"01111011", 
"10010001", 
"10000111", 
"10000000", 
"10010111", 
"01111011", 
"10001111", 
"01010100", 
"01101001", 
"01010010", 
"01101101", 
"10010101", 
"10000110", 
"10010011", 
"10110000", 
"01110101", 
"01111101", 
"10000111", 
"01101011", 
"01110001", 
"10001000", 
"01111011", 
"10010011", 
"01111000", 
"01111000", 
"00110001", 
"10011011", 
"10010001", 
"01111010", 
"10011101", 
"01010101", 
"01111110", 
"10011111", 
"01100101", 
"10000001", 
"10001000", 
"01000010", 
"01101110", 
"01111111", 
"10000001", 
"10000111", 
"10100100", 
"10001111", 
"10100111", 
"10000111", 
"10100000", 
"01011000", 
"10000001", 
"10010000", 
"01110101", 
"10010010", 
"01111011", 
"10000011", 
"01110010", 
"01111000", 
"10010000", 
"10000100", 
"10000101", 
"10001101", 
"10110101", 
"10010010", 
"10001111", 
"10001000", 
"10011000", 
"10100000", 
"10101110", 
"10001111", 
"01101000", 
"10010000", 
"01101101", 
"10001011", 
"10001000", 
"01100101", 
"10001101", 
"10000001", 
"00110110", 
"01111010", 
"10001010", 
"10010011", 
"10011110", 
"10001010", 
"10101011", 
"01111100", 
"01100101", 
"01010101", 
"01100011", 
"01101100", 
"01100100", 
"10000111", 
"01011010", 
"01110101", 
"01110111", 
"10001100", 
"01011111", 
"10001001", 
"01110111", 
"01100011", 
"00101010", 
"01110110", 
"10000110", 
"01111001", 
"01011111", 
"01110011", 
"10010000", 
"01110001", 
"10000010", 
"01000000", 
"01100010", 
"10010100", 
"01110001", 
"01111000", 
"01010000", 
"01101101", 
"01010101", 
"10001011", 
"01101110", 
"01111000", 
"01100101", 
"10000111", 
"10010000", 
"01111100", 
"01101100", 
"10010001", 
"10011110", 
"10010101", 
"01110101", 
"01111111", 
"01110101", 
"10010000", 
"10000011", 
"10000101", 
"01110100", 
"01011111", 
"10000100", 
"10000101", 
"10010111", 
"10000111", 
"10001000", 
"10001111", 
"01011111", 
"10001000", 
"01111001", 
"01100110", 
"10001011", 
"10000000", 
"01001100", 
"10001101", 
"10011111", 
"01011101", 
"10001111", 
"01110001", 
"10100111", 
"10001101", 
"10010010", 
"10001000", 
"10010101", 
"01111111", 
"10010111", 
"10000010", 
"10001001", 
"00111001", 
"00110100", 
"01111001", 
"10101010", 
"10101100", 
"01110100", 
"10000100", 
"01011110", 
"01101111", 
"10111110", 
"10001110", 
"10111111", 
"10001100", 
"01111011", 
"10101111", 
"10000100", 
"00001001", 
"00001111", 
"01111001", 
"01111011", 
"10011010", 
"01110011", 
"10000100", 
"01001001", 
"01110011", 
"10100111", 
"01011001", 
"01111110", 
"10001101", 
"10000000", 
"10011101", 
"01111010", 
"01001010", 
"00010010", 
"10000110", 
"10001001", 
"10001111", 
"10100000", 
"01110011", 
"01011101", 
"10001011", 
"01010000", 
"00111100", 
"01110111", 
"10000101", 
"01101100", 
"01111001", 
"01110011", 
"01010110", 
"01000111", 
"10010001", 
"01101110", 
"01010101", 
"10011001", 
"01111101", 
"01001111", 
"10110101", 
"00100111", 
"01100000", 
"10110010", 
"01110100", 
"10000011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_12: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_12(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
