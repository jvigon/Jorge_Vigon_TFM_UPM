use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_24_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_24_LAYER;

architecture Behavioral of ROM_FC_84_24_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_24: ROM_ARRAY_PESOS_FC_84 := (
"10100000", 
"00101111", 
"01011101", 
"10001011", 
"01101001", 
"10000011", 
"10011111", 
"01101110", 
"01011101", 
"10000010", 
"01100100", 
"01110101", 
"01111001", 
"01010010", 
"01100101", 
"01010101", 
"10001011", 
"01101111", 
"01111101", 
"01010100", 
"01110011", 
"01100111", 
"10000110", 
"01101101", 
"10000101", 
"10011010", 
"10000001", 
"10001110", 
"01110001", 
"01111100", 
"01011111", 
"01100111", 
"01111001", 
"01011010", 
"01100011", 
"01011011", 
"10000001", 
"01010010", 
"01100010", 
"10010000", 
"01100111", 
"01110111", 
"01110001", 
"01101101", 
"01011111", 
"10001101", 
"01101100", 
"10011000", 
"10000100", 
"10001011", 
"10011111", 
"10101010", 
"10010010", 
"01100001", 
"01101110", 
"10000101", 
"10010100", 
"01101110", 
"01011001", 
"10011011", 
"01101001", 
"00111001", 
"10001000", 
"01100100", 
"01111100", 
"01110111", 
"10010111", 
"01110011", 
"10010000", 
"10000010", 
"10010001", 
"01010110", 
"01100101", 
"01010111", 
"10001110", 
"01110110", 
"01001101", 
"10010101", 
"01101110", 
"01010001", 
"10000110", 
"01101010", 
"01111001", 
"01011011", 
"10001000", 
"10000010", 
"01100111", 
"10001000", 
"10000001", 
"10000110", 
"01001111", 
"01110100", 
"10010011", 
"01110111", 
"10000001", 
"01101001", 
"01000110", 
"10010011", 
"01101110", 
"10000110", 
"01100001", 
"10000011", 
"00101110", 
"01011000", 
"01111010", 
"01110001", 
"10001110", 
"01111001", 
"01011011", 
"01100111", 
"01100001", 
"01110001", 
"10000011", 
"01010110", 
"01100010", 
"10110101", 
"01101111", 
"10001001", 
"10000100", 
"01000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_24 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_24(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
