use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_67_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_67_LAYER;

architecture Behavioral of ROM_FC_120_67_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_67: ROM_ARRAY_PESOS_FC_120 := (
"01101100", 
"10000111", 
"01100101", 
"01100111", 
"01110001", 
"10000011", 
"01101001", 
"10000101", 
"01111100", 
"01111011", 
"01101101", 
"01111100", 
"01111010", 
"10001001", 
"01110101", 
"10000001", 
"10000000", 
"01101011", 
"01111010", 
"01110010", 
"01110011", 
"01110111", 
"01100110", 
"01110100", 
"01101011", 
"01111010", 
"10001101", 
"10000111", 
"01011001", 
"01110000", 
"10001000", 
"01111100", 
"01101011", 
"01111010", 
"01111001", 
"10000011", 
"10001110", 
"01101011", 
"01111101", 
"01111010", 
"01110010", 
"01110100", 
"01101000", 
"10000010", 
"10000010", 
"10000111", 
"01110010", 
"01101100", 
"01111010", 
"10000001", 
"01110001", 
"10000110", 
"01111101", 
"01110100", 
"01111100", 
"10000010", 
"10000101", 
"01011100", 
"01111010", 
"01101010", 
"10010101", 
"01110101", 
"01111011", 
"01101010", 
"01110111", 
"10000011", 
"10000001", 
"10001110", 
"10001110", 
"01111010", 
"10000011", 
"10001101", 
"10001100", 
"01100101", 
"10000001", 
"01110100", 
"01110010", 
"10001000", 
"10001010", 
"01111101", 
"01110001", 
"10001011", 
"01111011", 
"01100010", 
"01110111", 
"10000101", 
"01111011", 
"10001011", 
"01110010", 
"01111101", 
"01101010", 
"10001010", 
"01111010", 
"01111011", 
"10001100", 
"01110111", 
"01110000", 
"01101010", 
"01110111", 
"01111000", 
"01111010", 
"10000010", 
"01110111", 
"01111110", 
"10000110", 
"01110010", 
"10000001", 
"01101011", 
"01100100", 
"01100111", 
"01111100", 
"01111010", 
"10001111", 
"10000001", 
"01110000", 
"10001010", 
"10001101", 
"01110111", 
"01111011", 
"01100111", 
"01110011", 
"10001100", 
"01101111", 
"01110000", 
"01111110", 
"01110110", 
"01111000", 
"01110101", 
"10000111", 
"01110100", 
"10000011", 
"01101100", 
"10001110", 
"01111110", 
"10000011", 
"01101111", 
"01111011", 
"10001001", 
"10000110", 
"10001001", 
"01011110", 
"10000011", 
"01101010", 
"01101001", 
"10001010", 
"01111101", 
"01110011", 
"01101000", 
"10000110", 
"10000011", 
"10000001", 
"01110011", 
"10000011", 
"10001000", 
"01111011", 
"01110100", 
"10000011", 
"01111111", 
"01111100", 
"01110000", 
"01111111", 
"01101110", 
"01101001", 
"01100110", 
"01110111", 
"01111110", 
"10000100", 
"01101111", 
"10001011", 
"01110110", 
"10001010", 
"10000010", 
"01111010", 
"01101010", 
"01110101", 
"01101100", 
"10001100", 
"10000010", 
"01100111", 
"01110100", 
"01110011", 
"01101100", 
"10000010", 
"01111110", 
"01101001", 
"01110000", 
"01111110", 
"01101111", 
"01101101", 
"01110110", 
"01111110", 
"01111111", 
"10000001", 
"01111110", 
"10000000", 
"10101000", 
"01111100", 
"01110011", 
"01111111", 
"01101111", 
"10000001", 
"01110110", 
"01101000", 
"01111100", 
"01100101", 
"01111011", 
"01111101", 
"01110001", 
"01110101", 
"01101100", 
"01110101", 
"01101111", 
"10001010", 
"01101010", 
"01110111", 
"01101111", 
"10001111", 
"01110000", 
"10001000", 
"01111010", 
"01110011", 
"01111010", 
"10001001", 
"01111000", 
"01110100", 
"10001011", 
"01101001", 
"01100001", 
"10000111", 
"01101010", 
"10001100", 
"10000101", 
"01111010", 
"01100111", 
"01111110", 
"01101000", 
"01110010", 
"01110110", 
"10001001", 
"01101010", 
"10001101", 
"01010110", 
"10001110", 
"01110000", 
"10000001", 
"01100110", 
"01101111", 
"10000010", 
"10000110", 
"01111000", 
"01100110", 
"01110010", 
"01011111", 
"01110010", 
"10000010", 
"01110001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_67: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_67(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
