use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_35_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_35_LAYER;

architecture Behavioral of ROM_FC_84_35_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_35: ROM_ARRAY_PESOS_FC_84 := (
"01010110", 
"01000000", 
"10000011", 
"10001111", 
"10010100", 
"01111011", 
"01111011", 
"10001101", 
"10000000", 
"01001111", 
"10011011", 
"10010010", 
"01100101", 
"10000000", 
"10111010", 
"01100010", 
"01111000", 
"01100101", 
"01011110", 
"01000001", 
"10010011", 
"10010010", 
"10010000", 
"10010101", 
"01110110", 
"10011001", 
"01101111", 
"01100111", 
"10010110", 
"10010010", 
"10010000", 
"01010100", 
"01100101", 
"10100010", 
"01100011", 
"01110100", 
"01101110", 
"01101100", 
"10100100", 
"10000001", 
"01110111", 
"11100011", 
"01100011", 
"01110011", 
"10011111", 
"01010000", 
"10011100", 
"10010110", 
"01110101", 
"10101011", 
"01110101", 
"10101000", 
"01011001", 
"01100000", 
"10000100", 
"10011011", 
"11000011", 
"10011001", 
"01100010", 
"01111011", 
"01000101", 
"01011010", 
"10001001", 
"01101111", 
"01110101", 
"01011110", 
"10011100", 
"10000001", 
"01110011", 
"10001001", 
"01110100", 
"01110110", 
"01010001", 
"01001000", 
"10010011", 
"10001010", 
"01111110", 
"10101000", 
"10101011", 
"10010010", 
"01100111", 
"10010010", 
"10001000", 
"10010010", 
"01110111", 
"01110001", 
"01011010", 
"01100110", 
"10010011", 
"10010000", 
"10000101", 
"11101000", 
"01111010", 
"10010110", 
"01010010", 
"01111111", 
"01101010", 
"11010000", 
"01110001", 
"01110111", 
"10011001", 
"10000011", 
"10000100", 
"01011100", 
"10000011", 
"10010110", 
"01111011", 
"10010110", 
"01010000", 
"10101101", 
"01110011", 
"10001011", 
"10000110", 
"01110000", 
"01101100", 
"01110001", 
"01101101", 
"01011010", 
"01110111", 
"01011010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_35 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_35(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
