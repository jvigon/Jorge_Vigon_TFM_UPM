use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_32_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_32_LAYER;

architecture Behavioral of ROM_FC_120_32_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_32: ROM_ARRAY_PESOS_FC_120 := (
"01110101", 
"01010110", 
"01101101", 
"11000001", 
"01110110", 
"01110111", 
"10001011", 
"01110111", 
"01110101", 
"01110000", 
"01110010", 
"01100100", 
"01101110", 
"01110001", 
"10000111", 
"10001001", 
"01110111", 
"10010111", 
"10001010", 
"10100001", 
"01110011", 
"01101011", 
"10000011", 
"01111001", 
"01110001", 
"10001000", 
"10010000", 
"01010011", 
"01101010", 
"01110101", 
"01110011", 
"01110101", 
"10001001", 
"10000000", 
"01111011", 
"01100101", 
"10010000", 
"01011100", 
"01000100", 
"01110011", 
"01110001", 
"10001011", 
"10001011", 
"01110110", 
"01100110", 
"01100101", 
"01111101", 
"01101101", 
"01101001", 
"10000100", 
"01011111", 
"01011100", 
"01111100", 
"01011000", 
"00110011", 
"01110111", 
"10000010", 
"01110010", 
"01110011", 
"10010010", 
"01010010", 
"11000000", 
"01101111", 
"01110100", 
"01100100", 
"10001001", 
"01010101", 
"10001111", 
"01101010", 
"01100001", 
"10011110", 
"01111101", 
"01110011", 
"10001001", 
"01001101", 
"01011100", 
"10010100", 
"01100000", 
"10000010", 
"10001010", 
"01101101", 
"01000101", 
"01110011", 
"10100100", 
"10001011", 
"10001101", 
"01110000", 
"01111000", 
"10000111", 
"01110011", 
"01110000", 
"01001101", 
"10101011", 
"01101101", 
"10001010", 
"10000000", 
"01110010", 
"01001110", 
"01110001", 
"10001110", 
"10000000", 
"01111111", 
"10000010", 
"01110000", 
"10000010", 
"01111111", 
"01101011", 
"01011000", 
"01111000", 
"01001100", 
"01111011", 
"10000111", 
"10000010", 
"01001000", 
"01101110", 
"01001000", 
"01110011", 
"10000110", 
"01011110", 
"01011110", 
"01110110", 
"01011100", 
"01110000", 
"01110000", 
"01110111", 
"01001011", 
"01101011", 
"01110011", 
"01111001", 
"10001001", 
"01001100", 
"01110101", 
"10011000", 
"01101101", 
"10100001", 
"01110101", 
"10001001", 
"01111110", 
"10010111", 
"01100000", 
"10011010", 
"01000010", 
"01111011", 
"10001000", 
"01011100", 
"01101101", 
"01011001", 
"01101111", 
"10001111", 
"01111001", 
"01100110", 
"10001110", 
"01101101", 
"10101001", 
"10001110", 
"01111011", 
"01100111", 
"01001110", 
"10001001", 
"10000110", 
"01111010", 
"01011010", 
"01101101", 
"10001101", 
"10001011", 
"01101110", 
"01001010", 
"10000110", 
"10001110", 
"10001011", 
"01110011", 
"10010110", 
"01100110", 
"10001111", 
"01110010", 
"01110111", 
"01101100", 
"01110011", 
"10010111", 
"10010000", 
"10001010", 
"01010101", 
"01110010", 
"01111111", 
"10000101", 
"01101010", 
"10000100", 
"10100111", 
"10001000", 
"01011010", 
"01111111", 
"01111000", 
"10000101", 
"01001010", 
"01110011", 
"10111101", 
"01111101", 
"01110110", 
"01110000", 
"01101011", 
"10001011", 
"01101111", 
"10000010", 
"01010101", 
"00110100", 
"01011100", 
"01110011", 
"10000100", 
"10000101", 
"01100100", 
"01110110", 
"10110001", 
"10001100", 
"01111100", 
"01110100", 
"01111111", 
"01111111", 
"01110011", 
"01111011", 
"01100110", 
"10010000", 
"10001101", 
"10000110", 
"10000110", 
"01101011", 
"01011101", 
"01011011", 
"01010100", 
"10001101", 
"01101011", 
"01110100", 
"01111110", 
"01110000", 
"01110000", 
"01110001", 
"10001111", 
"10011100", 
"10001111", 
"10000110", 
"01110110", 
"01100110", 
"10001010", 
"01101011", 
"10100001", 
"01110110", 
"01110101", 
"01011001", 
"10000111", 
"01111011", 
"10001111", 
"10010100", 
"10001100", 
"10101111", 
"10000111", 
"10001100", 
"01110001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_32: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_32(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
