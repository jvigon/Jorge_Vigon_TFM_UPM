use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_45_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_45_LAYER;

architecture Behavioral of ROM_FC_120_45_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_45: ROM_ARRAY_PESOS_FC_120 := (
"01110111", 
"11000111", 
"01101011", 
"10110000", 
"10000000", 
"11101110", 
"10001001", 
"10001001", 
"01110010", 
"00110010", 
"01111010", 
"01010111", 
"01011100", 
"10101111", 
"01110001", 
"10011100", 
"10110100", 
"10010111", 
"01111000", 
"11001000", 
"01101100", 
"11000011", 
"10001110", 
"01001010", 
"10001111", 
"01101011", 
"01100000", 
"01100111", 
"01000100", 
"11111111", 
"10000010", 
"10000101", 
"10011110", 
"01110001", 
"01100000", 
"10101100", 
"01111001", 
"10011110", 
"11101010", 
"01110010", 
"01110101", 
"01000001", 
"01101011", 
"00111011", 
"00111001", 
"01101000", 
"10001110", 
"01101000", 
"10100110", 
"00111010", 
"10100010", 
"10001111", 
"10011000", 
"10100111", 
"11010011", 
"01111010", 
"10001001", 
"10101100", 
"01110111", 
"01111001", 
"01111111", 
"01101011", 
"01101010", 
"01101001", 
"01110000", 
"10000000", 
"10101101", 
"10000011", 
"10010100", 
"10011000", 
"01111110", 
"01110110", 
"01110010", 
"10010100", 
"10000001", 
"10001111", 
"11000000", 
"01111001", 
"01111111", 
"10100000", 
"01111011", 
"01110111", 
"10010100", 
"10010101", 
"01111000", 
"10001100", 
"10001000", 
"10000101", 
"10000100", 
"10101011", 
"10001010", 
"01110101", 
"10010000", 
"10000001", 
"01110100", 
"10001110", 
"01011111", 
"01001010", 
"10100011", 
"10110001", 
"01110111", 
"01101101", 
"10010100", 
"10001010", 
"10101101", 
"01001111", 
"01110111", 
"01011011", 
"01101011", 
"01100011", 
"01111111", 
"01011011", 
"10001000", 
"00101010", 
"01111010", 
"10100001", 
"01101101", 
"01111011", 
"10011011", 
"01110110", 
"10000001", 
"10011011", 
"10010000", 
"00110010", 
"00101110", 
"01110110", 
"01110110", 
"10000011", 
"01101111", 
"01110011", 
"10000010", 
"01110101", 
"10000111", 
"01111101", 
"01100001", 
"01101110", 
"01111001", 
"10110010", 
"10011010", 
"10000101", 
"01101100", 
"01100100", 
"10001110", 
"01111111", 
"01111111", 
"10011101", 
"10010010", 
"10010110", 
"10000011", 
"01111110", 
"01101010", 
"01101011", 
"01101111", 
"10001110", 
"10010111", 
"10100100", 
"01110001", 
"10101010", 
"10000010", 
"10001001", 
"10000110", 
"10010101", 
"10010001", 
"10001000", 
"01110100", 
"01110010", 
"10000110", 
"01001110", 
"10000111", 
"10100101", 
"01110100", 
"10000000", 
"10001111", 
"10110101", 
"01110011", 
"10010011", 
"01010100", 
"01000000", 
"01110101", 
"01101110", 
"01111100", 
"10011001", 
"01100011", 
"01110000", 
"10010000", 
"11000000", 
"10100011", 
"01011110", 
"10010001", 
"01000111", 
"01110111", 
"10010000", 
"01101100", 
"10110100", 
"00101000", 
"01100111", 
"10001100", 
"10000000", 
"10100101", 
"10100001", 
"10000111", 
"10011000", 
"10001011", 
"10001111", 
"10101000", 
"10011010", 
"01111111", 
"10000101", 
"10100011", 
"10011111", 
"01100101", 
"01101000", 
"01110100", 
"01101101", 
"01100010", 
"01011011", 
"01110101", 
"01100010", 
"01110011", 
"10100111", 
"01101110", 
"10000100", 
"10001101", 
"01111000", 
"10010111", 
"01111011", 
"01011010", 
"00110111", 
"10010010", 
"01110111", 
"01011001", 
"10010001", 
"10010010", 
"10001111", 
"10001001", 
"10001011", 
"01000100", 
"10011100", 
"01111101", 
"10001111", 
"01100000", 
"01001111", 
"01110100", 
"10000001", 
"10000101", 
"01110100", 
"01011110", 
"01111011", 
"01110010", 
"01110100", 
"10011011", 
"10010001", 
"01110111", 
"10110000", 
"10001010", 
"01111100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_45: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_45(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
