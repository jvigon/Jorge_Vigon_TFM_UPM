use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_111_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_111_LAYER;

architecture Behavioral of ROM_FC_120_111_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_111: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"10000000", 
"10000001", 
"10001011", 
"10001101", 
"10000011", 
"01101111", 
"10000111", 
"01111001", 
"10000101", 
"01100110", 
"01111111", 
"10011000", 
"10001100", 
"10001001", 
"10001110", 
"01101100", 
"01111001", 
"01100111", 
"01111011", 
"01101111", 
"01100100", 
"01111001", 
"10000011", 
"01101010", 
"01110011", 
"01111000", 
"01111010", 
"10000001", 
"01110010", 
"10001111", 
"01111101", 
"01110110", 
"01011010", 
"10001110", 
"10011000", 
"01101011", 
"01111111", 
"10000000", 
"10001010", 
"01101110", 
"01110001", 
"01101100", 
"01010010", 
"01111111", 
"01100111", 
"10000110", 
"01110101", 
"01111101", 
"01101010", 
"10001000", 
"01000001", 
"10001111", 
"01111001", 
"10000010", 
"01101100", 
"10001100", 
"01101110", 
"01101100", 
"10000011", 
"01111000", 
"01110100", 
"01110111", 
"10010001", 
"01101111", 
"01110101", 
"01110101", 
"01001110", 
"10001001", 
"01100111", 
"01100001", 
"01110001", 
"10001000", 
"01100110", 
"01111101", 
"10001001", 
"01110100", 
"01110110", 
"01111010", 
"01111011", 
"01111110", 
"01110110", 
"01110111", 
"01000110", 
"10000110", 
"01110110", 
"01101011", 
"01100111", 
"01111001", 
"01111000", 
"10000010", 
"01111101", 
"01101010", 
"01011101", 
"01111010", 
"01101010", 
"01110110", 
"10001001", 
"10001001", 
"01110001", 
"01101011", 
"01111010", 
"01110001", 
"10000100", 
"01110010", 
"01100011", 
"01111001", 
"01101110", 
"01100000", 
"01101101", 
"10001101", 
"10000101", 
"01100110", 
"10000101", 
"10000111", 
"01001010", 
"01111001", 
"01011101", 
"01111110", 
"10000111", 
"01111000", 
"01100001", 
"01110100", 
"01111110", 
"01110111", 
"10010100", 
"10001110", 
"01110101", 
"01110100", 
"10001010", 
"01100000", 
"01100001", 
"10000001", 
"10010100", 
"01101101", 
"01101001", 
"10000101", 
"01100111", 
"10000101", 
"10001011", 
"01011111", 
"10000010", 
"10001011", 
"01110011", 
"01111000", 
"10000001", 
"10000000", 
"01110010", 
"10010000", 
"01110111", 
"01101011", 
"01111110", 
"01110110", 
"01010010", 
"10001110", 
"01110010", 
"01100011", 
"01111000", 
"10001011", 
"10001010", 
"01101001", 
"10000111", 
"10001101", 
"10001101", 
"01101101", 
"01110110", 
"10000101", 
"01111000", 
"01110010", 
"01101011", 
"01110011", 
"10000001", 
"10000010", 
"10000111", 
"01111111", 
"01111001", 
"01101100", 
"01111100", 
"01101110", 
"10011000", 
"10001000", 
"01101101", 
"10001001", 
"10000100", 
"01110000", 
"01101011", 
"01100111", 
"01110111", 
"01101000", 
"10000110", 
"10001000", 
"10001100", 
"01110011", 
"01100100", 
"01100101", 
"00101111", 
"01111001", 
"10000000", 
"01101110", 
"10000110", 
"01101010", 
"10001000", 
"10010001", 
"01100010", 
"01011101", 
"01101010", 
"01111001", 
"01110100", 
"10001011", 
"01100100", 
"10000100", 
"01111101", 
"10000101", 
"01110101", 
"01011001", 
"01101101", 
"01110010", 
"01110010", 
"01110111", 
"01100101", 
"10000000", 
"10001010", 
"10000001", 
"10001011", 
"01110001", 
"01110111", 
"01110010", 
"01110001", 
"01110001", 
"10000011", 
"01101010", 
"10000111", 
"10001011", 
"10000101", 
"01101111", 
"01110101", 
"00111100", 
"01110000", 
"01110111", 
"01111011", 
"01101001", 
"01101000", 
"01111111", 
"10001010", 
"10001011", 
"01101110", 
"01101101", 
"01110000", 
"10001011", 
"01111100", 
"01110111", 
"11000001", 
"01100010", 
"10000000", 
"01110100", 
"01111000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_111 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_111(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
