use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_85_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_85_LAYER;

architecture Behavioral of ROM_FC_120_85_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_85: ROM_ARRAY_PESOS_FC_120 := (
"01101101", 
"01110100", 
"11001001", 
"10100100", 
"01110100", 
"01111010", 
"01101100", 
"01101101", 
"10000110", 
"10011000", 
"01101001", 
"01011011", 
"01111110", 
"10100100", 
"10011001", 
"10000001", 
"10000101", 
"01111100", 
"01101001", 
"01010111", 
"01111100", 
"01110010", 
"01111011", 
"01101000", 
"01111001", 
"10000100", 
"01011011", 
"01101100", 
"10010011", 
"10011010", 
"10010000", 
"01111100", 
"10000110", 
"01001100", 
"10000010", 
"10010111", 
"01101101", 
"01110001", 
"01100111", 
"01111011", 
"01110110", 
"01110100", 
"01111011", 
"01100001", 
"10001011", 
"10010100", 
"01110111", 
"10010001", 
"01110111", 
"01110011", 
"10001111", 
"01110010", 
"01111010", 
"10001110", 
"01001110", 
"10000010", 
"10010011", 
"01001011", 
"01110011", 
"01110000", 
"10000110", 
"10010111", 
"01111001", 
"01111101", 
"10000001", 
"10010011", 
"01101010", 
"00111110", 
"10000001", 
"01111101", 
"10000111", 
"10000001", 
"10000101", 
"10011000", 
"10011111", 
"01101100", 
"10000101", 
"01001110", 
"10010011", 
"10010011", 
"10001010", 
"10010010", 
"01100110", 
"00111010", 
"01101111", 
"01111100", 
"01111110", 
"10000001", 
"01110100", 
"10010001", 
"10110000", 
"10001001", 
"01010111", 
"01101111", 
"10000010", 
"10001101", 
"01110010", 
"10010000", 
"01111011", 
"01101110", 
"01111100", 
"01101011", 
"01110011", 
"01111010", 
"10000011", 
"10001100", 
"01111111", 
"01011101", 
"10000011", 
"01101100", 
"01111111", 
"10000101", 
"01100001", 
"10011111", 
"01100101", 
"10100001", 
"01111110", 
"10000001", 
"01010001", 
"10000001", 
"01101110", 
"01110100", 
"10001011", 
"01111100", 
"01110110", 
"10011011", 
"10001101", 
"10010101", 
"01110100", 
"01011111", 
"01100001", 
"01001000", 
"10001111", 
"10010010", 
"10000111", 
"10100001", 
"10001111", 
"01101001", 
"01100111", 
"01100100", 
"10010101", 
"10010100", 
"10000100", 
"01101101", 
"10001001", 
"10001000", 
"01110110", 
"01010110", 
"10000111", 
"10001100", 
"10001111", 
"10011101", 
"01101110", 
"01010001", 
"01101011", 
"10000101", 
"10001101", 
"10001111", 
"01111101", 
"10010101", 
"01101001", 
"01110100", 
"10001111", 
"01110111", 
"01111001", 
"10010011", 
"10100101", 
"01100011", 
"10001111", 
"01111000", 
"01100110", 
"10001000", 
"10001101", 
"01110010", 
"01111001", 
"01111001", 
"10010011", 
"01101100", 
"01101101", 
"01110111", 
"01110111", 
"10000001", 
"01101111", 
"01010100", 
"10001110", 
"10000101", 
"10001100", 
"01011110", 
"10111110", 
"01101010", 
"10000110", 
"01111010", 
"10000001", 
"01110110", 
"01101000", 
"01010110", 
"01110101", 
"10010001", 
"01110111", 
"10011100", 
"01110110", 
"10001000", 
"01110011", 
"01010011", 
"01010110", 
"10000100", 
"01110000", 
"01111001", 
"01110111", 
"10000110", 
"01100001", 
"01111000", 
"10000001", 
"10010011", 
"10001001", 
"01100011", 
"10001001", 
"01101111", 
"10010001", 
"01011100", 
"01011110", 
"01111101", 
"10001000", 
"10010011", 
"10010010", 
"01011011", 
"01110101", 
"01100110", 
"01110100", 
"10011110", 
"10010011", 
"01101100", 
"10000010", 
"01101011", 
"10000000", 
"01001011", 
"01010110", 
"01101011", 
"10010100", 
"01110001", 
"10000101", 
"01010001", 
"01100111", 
"01101111", 
"01110111", 
"01101100", 
"01011000", 
"10001111", 
"01110011", 
"10000001", 
"10101111", 
"10001000", 
"01001011", 
"01011010", 
"10000101", 
"01110100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_85: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_85(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
