use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_40_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_40_LAYER;

architecture Behavioral of ROM_FC_120_40_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_40: ROM_ARRAY_PESOS_FC_120 := (
"10000100", 
"01001011", 
"10011010", 
"10011111", 
"10011001", 
"00101110", 
"10000010", 
"10010001", 
"01111101", 
"10100000", 
"10101001", 
"01111111", 
"10101100", 
"10010001", 
"01111000", 
"10001110", 
"01111110", 
"01011010", 
"10000111", 
"10001101", 
"01100100", 
"00001011", 
"01100011", 
"10000111", 
"10001011", 
"10011001", 
"10000000", 
"01110101", 
"10010001", 
"01110101", 
"10001111", 
"10101001", 
"10000011", 
"01101100", 
"10011110", 
"01110010", 
"01110111", 
"01011100", 
"01001110", 
"10000010", 
"01110100", 
"01111110", 
"01010000", 
"01111010", 
"01111100", 
"10101110", 
"10000000", 
"10010100", 
"01101111", 
"10000010", 
"01010000", 
"00111110", 
"01110111", 
"01001111", 
"00111110", 
"01111000", 
"10001010", 
"10100100", 
"01001110", 
"01110000", 
"01110011", 
"10010010", 
"10000011", 
"01111111", 
"01110101", 
"10100101", 
"10111011", 
"10111010", 
"10000001", 
"10010110", 
"01101000", 
"01110001", 
"10000110", 
"10011000", 
"10001101", 
"00110110", 
"01101011", 
"01101000", 
"01110011", 
"10001010", 
"01011111", 
"10001010", 
"10000100", 
"01111110", 
"01100111", 
"10011001", 
"01110101", 
"10001011", 
"01111110", 
"10011010", 
"01110111", 
"01110000", 
"01111101", 
"11010000", 
"01101101", 
"10010001", 
"01101000", 
"10101110", 
"00110000", 
"00100011", 
"01111011", 
"01110110", 
"01110100", 
"01101100", 
"01100100", 
"10000111", 
"10001111", 
"10101001", 
"01111111", 
"10001111", 
"10100001", 
"10100101", 
"01111001", 
"01101111", 
"01001110", 
"01110011", 
"01110011", 
"10011101", 
"01111011", 
"10000110", 
"10000001", 
"01010010", 
"10010000", 
"10001101", 
"10011000", 
"10110001", 
"10010011", 
"01111110", 
"01110100", 
"01110000", 
"10011001", 
"01111010", 
"01100010", 
"01111101", 
"00111010", 
"01111000", 
"01101000", 
"01111001", 
"01110100", 
"10000100", 
"10000110", 
"01000001", 
"10001110", 
"01110001", 
"10010000", 
"01110001", 
"10100110", 
"10001111", 
"10000101", 
"10011100", 
"10001010", 
"10011101", 
"01100110", 
"10000001", 
"01111110", 
"10010000", 
"10001110", 
"10000110", 
"01101000", 
"10001100", 
"01101101", 
"01110010", 
"01110001", 
"01011001", 
"01110001", 
"10011111", 
"01110110", 
"01111101", 
"10000110", 
"01100010", 
"01001000", 
"01101100", 
"10001011", 
"01000010", 
"01110101", 
"10010001", 
"01110100", 
"01111111", 
"01010111", 
"10000111", 
"10000111", 
"10100010", 
"10000111", 
"01010100", 
"10010010", 
"01111010", 
"10001101", 
"01111110", 
"10011111", 
"01101111", 
"01101010", 
"10001101", 
"01100111", 
"01100001", 
"01000111", 
"00010110", 
"10000111", 
"01110101", 
"10000111", 
"10101011", 
"01111100", 
"10010000", 
"01110011", 
"10000011", 
"01100001", 
"01011101", 
"01110111", 
"10000101", 
"10001010", 
"01101100", 
"01101001", 
"00101110", 
"10001100", 
"10100110", 
"10001001", 
"10010000", 
"10011000", 
"01111110", 
"01110011", 
"01111101", 
"01101100", 
"01111010", 
"10001100", 
"01100101", 
"10010110", 
"01110001", 
"01101000", 
"01000101", 
"10100011", 
"10001110", 
"10001111", 
"10000110", 
"10110010", 
"10010100", 
"01010001", 
"10100000", 
"10000100", 
"10010100", 
"10001010", 
"01110011", 
"01011001", 
"01001001", 
"10000011", 
"01100111", 
"10000100", 
"10000000", 
"10010101", 
"01110110", 
"10010111", 
"01011111", 
"10100000", 
"01111111", 
"00111111", 
"00110010", 
"01111010", 
"10000011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_40: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_40(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
