use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_26_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_26_LAYER;

architecture Behavioral of ROM_FC_120_26_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_26: ROM_ARRAY_PESOS_FC_120 := (
"01110010", 
"01110011", 
"01100100", 
"10110100", 
"01111110", 
"01110100", 
"10011111", 
"01011110", 
"10000100", 
"10010111", 
"01110101", 
"01011001", 
"10010100", 
"10000101", 
"10010001", 
"01101100", 
"10011010", 
"01111101", 
"10010000", 
"10001100", 
"10010001", 
"11000001", 
"01001100", 
"01010010", 
"01101111", 
"10000011", 
"01110101", 
"10101011", 
"10000010", 
"11000010", 
"01111001", 
"10000011", 
"01110011", 
"01111101", 
"10001001", 
"10000000", 
"01101011", 
"01000010", 
"10000001", 
"01011110", 
"10001000", 
"10001001", 
"01001110", 
"10010100", 
"01111000", 
"10011111", 
"01110110", 
"01110010", 
"01110111", 
"01111100", 
"01101100", 
"10010010", 
"01110110", 
"01111001", 
"01110110", 
"01111010", 
"10000010", 
"10001000", 
"01101101", 
"10111101", 
"01110010", 
"10101111", 
"01111011", 
"01100011", 
"01010111", 
"01100100", 
"10000100", 
"01100011", 
"10100010", 
"10001000", 
"10000111", 
"00110010", 
"10010100", 
"01111000", 
"01110100", 
"01100001", 
"10100110", 
"10000101", 
"10010111", 
"10011110", 
"01110011", 
"10001110", 
"01111100", 
"10010001", 
"01111001", 
"01010100", 
"10001100", 
"01101011", 
"01110101", 
"10001010", 
"10011111", 
"10001011", 
"10010100", 
"10011101", 
"10001110", 
"01111011", 
"10010000", 
"10001011", 
"10011001", 
"10101000", 
"10001000", 
"01101011", 
"10010010", 
"01110111", 
"01111001", 
"10001011", 
"01001011", 
"01111110", 
"10011111", 
"01111001", 
"10000110", 
"10001011", 
"10011111", 
"10001000", 
"01100000", 
"01001011", 
"10001010", 
"01100010", 
"01010011", 
"10000111", 
"01111011", 
"10011101", 
"01001111", 
"01100010", 
"10010111", 
"01100101", 
"01111111", 
"10010011", 
"10000000", 
"10000011", 
"01011011", 
"01100010", 
"01110000", 
"01100110", 
"01011110", 
"01101100", 
"01010111", 
"01111010", 
"10001001", 
"01111011", 
"10001111", 
"01110011", 
"10001111", 
"10011000", 
"01011010", 
"01011001", 
"01110101", 
"01110111", 
"01110101", 
"01100110", 
"10010001", 
"10101001", 
"10010010", 
"01101011", 
"01101111", 
"01001110", 
"10010001", 
"01101000", 
"10001100", 
"01110010", 
"10011110", 
"00110111", 
"10000111", 
"10011000", 
"10000000", 
"10010010", 
"01010111", 
"01100011", 
"01101100", 
"01111111", 
"10001001", 
"10011000", 
"01111100", 
"11100001", 
"10000011", 
"10000010", 
"01111010", 
"10000001", 
"10000101", 
"01100110", 
"10001000", 
"01011101", 
"01011100", 
"10010100", 
"10000000", 
"10100000", 
"01010000", 
"01111010", 
"01100000", 
"01011110", 
"10001111", 
"01101101", 
"01011011", 
"11000001", 
"10011000", 
"01001000", 
"10001101", 
"01011100", 
"10011001", 
"01101110", 
"10001000", 
"01011010", 
"01101101", 
"10001011", 
"10101100", 
"01101101", 
"10001101", 
"01101001", 
"01100100", 
"10110011", 
"10010100", 
"10001100", 
"10000111", 
"10001000", 
"10011110", 
"01100000", 
"01111111", 
"01011001", 
"01101010", 
"00111101", 
"10101001", 
"10001001", 
"10010010", 
"01111011", 
"01110100", 
"10001101", 
"01100110", 
"01011110", 
"01110111", 
"10000101", 
"01111100", 
"01100000", 
"10001001", 
"01100101", 
"10111001", 
"01100101", 
"10011110", 
"10100100", 
"10000101", 
"10000000", 
"01010111", 
"01111111", 
"01101100", 
"01110101", 
"10010100", 
"01110010", 
"10100001", 
"01101101", 
"01111001", 
"01000101", 
"01101010", 
"10001010", 
"01111101", 
"10011011", 
"01110011", 
"10001010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_26: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_26(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
