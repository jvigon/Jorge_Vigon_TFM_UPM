use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_102_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_102_LAYER;

architecture Behavioral of ROM_FC_120_102_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_102: ROM_ARRAY_PESOS_FC_120 := (
"01101001", 
"01010001", 
"01111010", 
"01100000", 
"10011000", 
"00100111", 
"10010011", 
"10010000", 
"01011101", 
"10010101", 
"10100001", 
"01111110", 
"10101101", 
"00100100", 
"10010010", 
"01111111", 
"00101111", 
"10000001", 
"10010111", 
"10110111", 
"10001111", 
"00000000", 
"10001110", 
"10000100", 
"01101110", 
"10001101", 
"10010001", 
"10110011", 
"10011100", 
"00000000", 
"01111000", 
"10010001", 
"01100000", 
"10010001", 
"10011101", 
"10000101", 
"01110100", 
"01101000", 
"01011110", 
"10000110", 
"01110000", 
"01110101", 
"01100010", 
"10000010", 
"10100010", 
"01110001", 
"01111101", 
"01110010", 
"10000111", 
"10101001", 
"00101100", 
"01010110", 
"01010101", 
"01010000", 
"01000011", 
"10010101", 
"01110000", 
"01101000", 
"01100011", 
"00010100", 
"01100101", 
"10100101", 
"01101000", 
"01010100", 
"10000000", 
"00011110", 
"10001000", 
"10100000", 
"10001011", 
"10010001", 
"01110010", 
"10011100", 
"01011010", 
"01110101", 
"01111101", 
"00000011", 
"00000000", 
"10010101", 
"01011010", 
"10001111", 
"00101111", 
"01101010", 
"10010000", 
"10100010", 
"10001101", 
"10000001", 
"10010111", 
"01100011", 
"01111101", 
"01101110", 
"01111010", 
"10000010", 
"01111011", 
"11000100", 
"10001111", 
"01110001", 
"01100001", 
"10100110", 
"10010010", 
"01111011", 
"01111111", 
"10110100", 
"10011011", 
"10100001", 
"01111011", 
"01110001", 
"10010100", 
"10000110", 
"10011000", 
"01100001", 
"01110101", 
"01110000", 
"10010000", 
"10100011", 
"01101110", 
"01101100", 
"10001000", 
"10100011", 
"11010010", 
"10110101", 
"10001011", 
"00111000", 
"01111011", 
"01001011", 
"10001110", 
"01101000", 
"10000110", 
"01110110", 
"10011000", 
"01101110", 
"10010111", 
"10010100", 
"01001001", 
"01011010", 
"01010111", 
"01001101", 
"10001101", 
"01110011", 
"01000101", 
"01010000", 
"01010100", 
"10110010", 
"10010010", 
"01111000", 
"01000110", 
"01101010", 
"10000101", 
"10000001", 
"10000101", 
"01101011", 
"01101111", 
"01011001", 
"10000010", 
"10110011", 
"01101010", 
"10010010", 
"10001101", 
"10001111", 
"01110111", 
"01110100", 
"01001101", 
"10000100", 
"10001101", 
"01111100", 
"01110101", 
"10110100", 
"01101101", 
"10011001", 
"10000000", 
"10010111", 
"01100111", 
"01011010", 
"10000100", 
"00110101", 
"10011111", 
"10010000", 
"10000010", 
"01111001", 
"01100001", 
"01111001", 
"01110000", 
"10101111", 
"10010011", 
"01111101", 
"01101011", 
"01010011", 
"10001011", 
"01000001", 
"01010101", 
"01101001", 
"10011010", 
"01110100", 
"01101101", 
"01110011", 
"01101111", 
"01110010", 
"01010010", 
"01010100", 
"10010010", 
"10001011", 
"10001100", 
"10000000", 
"10000101", 
"01111001", 
"10110101", 
"10000100", 
"01110001", 
"10001111", 
"10001110", 
"01100101", 
"00111101", 
"01000101", 
"01011111", 
"10010100", 
"10101100", 
"10001100", 
"01001111", 
"10011111", 
"01001110", 
"10011110", 
"10010010", 
"10001101", 
"01101110", 
"01110001", 
"10010111", 
"01110100", 
"01000000", 
"01011100", 
"01011110", 
"01111000", 
"01101111", 
"01101111", 
"10010010", 
"01010010", 
"01110010", 
"01110111", 
"01110000", 
"01010000", 
"10001001", 
"01111110", 
"10000011", 
"00101000", 
"10010100", 
"01011000", 
"10001100", 
"10001101", 
"10110000", 
"01111011", 
"01111110", 
"01001110", 
"01111000", 
"00110001", 
"00000000", 
"01010001", 
"01110000", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_102: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_102(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
