use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_5_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_5_LAYER;

architecture Behavioral of ROM_FC_120_5_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_5: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"10100010", 
"01111001", 
"10010000", 
"01111100", 
"01110110", 
"10100010", 
"10000010", 
"10001111", 
"01010110", 
"01111101", 
"01110010", 
"01101011", 
"01111101", 
"10001101", 
"10011100", 
"10100001", 
"01110010", 
"01110000", 
"10001000", 
"01100111", 
"10010001", 
"01100000", 
"10001101", 
"01111110", 
"01110111", 
"01101110", 
"01111001", 
"10010001", 
"10000100", 
"10010001", 
"10011101", 
"10100000", 
"01111100", 
"01100110", 
"01100010", 
"01101011", 
"01011011", 
"01101000", 
"10000110", 
"10001010", 
"01011110", 
"01101110", 
"10011011", 
"10000010", 
"01101110", 
"01110011", 
"01100100", 
"10000100", 
"01001110", 
"10010101", 
"01010011", 
"10000101", 
"01110100", 
"10010010", 
"01111010", 
"10000100", 
"10001110", 
"01101111", 
"10000100", 
"10001000", 
"01111010", 
"01111000", 
"10000010", 
"10001001", 
"01110010", 
"01110111", 
"01101110", 
"10000100", 
"01011001", 
"10010001", 
"01100100", 
"01111000", 
"10001101", 
"01101001", 
"01001011", 
"10100001", 
"01111110", 
"01110010", 
"10001000", 
"01100011", 
"10000011", 
"01111000", 
"01010011", 
"01111110", 
"10101010", 
"01110011", 
"10000110", 
"01111110", 
"01101011", 
"01110001", 
"01001101", 
"10001110", 
"01101011", 
"01111000", 
"10000000", 
"01100101", 
"01110100", 
"10001011", 
"01000011", 
"01110111", 
"01110110", 
"01101100", 
"01100010", 
"01111000", 
"10010000", 
"10010000", 
"01100101", 
"01110101", 
"01111100", 
"01101111", 
"01110101", 
"01111110", 
"10100001", 
"01111101", 
"00111111", 
"01111010", 
"01101101", 
"10000111", 
"01001110", 
"10010010", 
"10110111", 
"10000000", 
"10001111", 
"11000010", 
"01011111", 
"01101101", 
"10000000", 
"10000110", 
"10001000", 
"01110111", 
"01011111", 
"01110010", 
"10001110", 
"10010101", 
"01110001", 
"01110111", 
"01110101", 
"01100100", 
"10000011", 
"10000011", 
"01011111", 
"01111110", 
"10000111", 
"01110100", 
"10001101", 
"01100111", 
"01000110", 
"10000001", 
"10001110", 
"01100110", 
"10001000", 
"01111011", 
"01100110", 
"01110110", 
"10000100", 
"01110100", 
"01101110", 
"10010001", 
"10000010", 
"10001001", 
"10001100", 
"01111110", 
"01100011", 
"01101010", 
"10001010", 
"10000000", 
"10001000", 
"01101110", 
"01101001", 
"01110101", 
"01101001", 
"10000111", 
"10001001", 
"01111111", 
"01101001", 
"01101010", 
"10001011", 
"01110101", 
"01101100", 
"10000001", 
"10000000", 
"01100101", 
"10000100", 
"10000011", 
"01011000", 
"01110100", 
"10000110", 
"10000001", 
"10000010", 
"01101000", 
"01111000", 
"10001000", 
"01111011", 
"01101011", 
"01010010", 
"10010001", 
"10010000", 
"01101110", 
"01101011", 
"01111100", 
"10010101", 
"01111000", 
"01010111", 
"10100111", 
"10011000", 
"01110111", 
"10001000", 
"10000101", 
"01110011", 
"01111111", 
"01011000", 
"10001011", 
"10010100", 
"10000100", 
"10011100", 
"10001010", 
"10001100", 
"01110010", 
"01010101", 
"10000001", 
"10001111", 
"01111001", 
"10001111", 
"10000110", 
"01001111", 
"01101001", 
"01011100", 
"01111110", 
"01100111", 
"10001010", 
"01111011", 
"01101100", 
"01101110", 
"01110011", 
"01011011", 
"10000100", 
"01110100", 
"10000101", 
"01110010", 
"10000110", 
"01001100", 
"10000000", 
"01110110", 
"01111010", 
"01110111", 
"01011000", 
"10010010", 
"10000111", 
"01011011", 
"01110001", 
"01111100", 
"01101101", 
"01110100", 
"10000010", 
"01111001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_5 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_5(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
