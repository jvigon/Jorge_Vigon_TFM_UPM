use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_95_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_95_LAYER;

architecture Behavioral of ROM_FC_120_95_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_95: ROM_ARRAY_PESOS_FC_120 := (
"01101000", 
"10000100", 
"01011100", 
"01100110", 
"10000101", 
"01111000", 
"01111101", 
"01100001", 
"01101101", 
"10000110", 
"01111101", 
"01101100", 
"01100111", 
"01111101", 
"10000000", 
"01111100", 
"01110100", 
"01100001", 
"01000011", 
"01101110", 
"01010111", 
"10000101", 
"10000100", 
"01110000", 
"10000000", 
"01011110", 
"01010010", 
"01110111", 
"01111001", 
"10000000", 
"10000101", 
"01110111", 
"01111000", 
"01110010", 
"01101001", 
"01110100", 
"01110001", 
"01110111", 
"01111001", 
"01101111", 
"10000101", 
"01101101", 
"01011100", 
"10001100", 
"01110100", 
"10000100", 
"10000110", 
"10010011", 
"01100011", 
"01010000", 
"01110011", 
"01111100", 
"10000100", 
"01001111", 
"10101001", 
"10000101", 
"01110110", 
"01110011", 
"01110111", 
"10000000", 
"10001110", 
"01000001", 
"10001101", 
"10001111", 
"01101011", 
"01010111", 
"01110010", 
"01111100", 
"10000001", 
"10011001", 
"01100110", 
"01111010", 
"10001011", 
"10001010", 
"01011101", 
"10000011", 
"01111011", 
"01111101", 
"10001001", 
"10000010", 
"01101000", 
"01110111", 
"01111110", 
"01110111", 
"01101000", 
"01110011", 
"01111110", 
"01110110", 
"01101010", 
"01101000", 
"01011101", 
"01100100", 
"01100100", 
"10001010", 
"01110010", 
"10001011", 
"01111011", 
"01011111", 
"01110000", 
"10000000", 
"01101101", 
"01100010", 
"10000111", 
"10001010", 
"01101011", 
"01111010", 
"01100100", 
"01111001", 
"01011111", 
"01101111", 
"10001101", 
"01110010", 
"01110101", 
"01100011", 
"01111101", 
"10001000", 
"10000011", 
"01110101", 
"01111101", 
"01101010", 
"01110111", 
"10110110", 
"01101001", 
"01111001", 
"01101011", 
"01101101", 
"01111000", 
"10001100", 
"10000011", 
"01100010", 
"01011101", 
"01110000", 
"10000010", 
"10000010", 
"01110010", 
"01111000", 
"10001111", 
"10001011", 
"01111111", 
"10000101", 
"01110110", 
"01101100", 
"10000110", 
"01101110", 
"10001100", 
"01110101", 
"01110011", 
"01111111", 
"01110100", 
"10010111", 
"01010101", 
"10001010", 
"01101001", 
"01100100", 
"01110010", 
"01111001", 
"01010110", 
"01111000", 
"01110111", 
"10000101", 
"10000111", 
"01110101", 
"01110100", 
"10000111", 
"10001001", 
"01011001", 
"01100010", 
"01111010", 
"01101000", 
"10010010", 
"01110011", 
"01101101", 
"01110111", 
"01100111", 
"10000100", 
"10001110", 
"01101111", 
"01100011", 
"01101110", 
"10000111", 
"01111011", 
"01011011", 
"10001000", 
"01111010", 
"10000001", 
"10001011", 
"01100111", 
"01101110", 
"10000000", 
"01110000", 
"01101110", 
"10001110", 
"01111110", 
"10000101", 
"01111110", 
"10000110", 
"01111000", 
"01111111", 
"01110000", 
"01100111", 
"01011111", 
"01101111", 
"01110011", 
"10011001", 
"10001101", 
"01110011", 
"01111011", 
"01111001", 
"01101010", 
"01110011", 
"01111110", 
"10000001", 
"10000010", 
"10000000", 
"01111000", 
"10011011", 
"10000000", 
"01110111", 
"10001000", 
"01101101", 
"01101101", 
"01011001", 
"10001011", 
"01101111", 
"01110000", 
"01100110", 
"01100000", 
"01110110", 
"10000111", 
"01001101", 
"01011100", 
"01101111", 
"01111010", 
"01110111", 
"01111101", 
"01011011", 
"01101101", 
"01111010", 
"01110100", 
"10000101", 
"01110010", 
"01011011", 
"01110101", 
"01110101", 
"01111101", 
"01101101", 
"01100001", 
"01100010", 
"10001010", 
"01011011", 
"01011111", 
"01111000", 
"10000011", 
"01101100", 
"01110001", 
"01110100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_95: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_95(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
