use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_20_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_20_LAYER;

architecture Behavioral of ROM_FC_84_20_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_20: ROM_ARRAY_PESOS_FC_84 := (
"01101000", 
"01110011", 
"10001011", 
"10001000", 
"01010100", 
"10011010", 
"10000111", 
"01111101", 
"10001000", 
"10011001", 
"10001001", 
"01001100", 
"01110101", 
"10110011", 
"10101000", 
"01110000", 
"00111101", 
"10000001", 
"10001001", 
"00110000", 
"10001111", 
"01100001", 
"01110110", 
"01001111", 
"10001100", 
"10111100", 
"10001000", 
"01010000", 
"01100110", 
"10010000", 
"01101101", 
"01110010", 
"10000000", 
"01111111", 
"01110000", 
"10001001", 
"01011110", 
"01101100", 
"01110101", 
"10010100", 
"01101001", 
"01100001", 
"01010110", 
"01001111", 
"10101111", 
"01101000", 
"10001011", 
"01111000", 
"01010111", 
"10010111", 
"01100100", 
"01110011", 
"01101100", 
"10010101", 
"01001011", 
"10101110", 
"10010011", 
"01101110", 
"01011000", 
"01000100", 
"01101110", 
"01110110", 
"10011011", 
"01001011", 
"10011110", 
"10001101", 
"11011100", 
"01100000", 
"01100111", 
"01110111", 
"00111110", 
"01001001", 
"10001000", 
"01011101", 
"01110001", 
"10011100", 
"01111100", 
"01111000", 
"01100111", 
"00111101", 
"01010010", 
"01100001", 
"01001001", 
"01000000", 
"01000000", 
"01101100", 
"01101010", 
"01111000", 
"01110111", 
"01001010", 
"01101011", 
"01101011", 
"10011000", 
"01101011", 
"01111100", 
"10000101", 
"01011010", 
"10000111", 
"10101000", 
"10001010", 
"10001010", 
"01110000", 
"01100111", 
"01100001", 
"01110111", 
"01111101", 
"00111110", 
"10010010", 
"01011111", 
"10000101", 
"10110110", 
"10010110", 
"10001000", 
"01100101", 
"01111001", 
"01011101", 
"10000101", 
"10001001", 
"10001000", 
"01110010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_20 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_20(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
