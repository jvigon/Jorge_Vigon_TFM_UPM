use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_45_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_45_LAYER;

architecture Behavioral of ROM_FC_84_45_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_45: ROM_ARRAY_PESOS_FC_84 := (
"10000001", 
"10010110", 
"10010010", 
"01111101", 
"10001111", 
"01101000", 
"10010111", 
"10000011", 
"01111000", 
"10100001", 
"01110000", 
"01100000", 
"10010101", 
"10000101", 
"01010001", 
"01011111", 
"01111101", 
"01101110", 
"00111111", 
"01010111", 
"10001111", 
"01010001", 
"10000111", 
"10000000", 
"01111011", 
"10011001", 
"10011010", 
"01011101", 
"01110110", 
"01110000", 
"10001011", 
"01101101", 
"01100111", 
"10000111", 
"10101101", 
"01001000", 
"10010011", 
"01111010", 
"01110011", 
"10010011", 
"01011111", 
"01101001", 
"01011110", 
"01111010", 
"01101001", 
"01101101", 
"01110000", 
"01101100", 
"01110111", 
"01111011", 
"01111100", 
"10001100", 
"10010011", 
"10000000", 
"01111111", 
"01110001", 
"10010011", 
"10000010", 
"01100000", 
"01111111", 
"01100001", 
"01001111", 
"10011000", 
"10011110", 
"01100110", 
"10010001", 
"01110110", 
"10000010", 
"01110001", 
"00110010", 
"01110010", 
"01010000", 
"00101000", 
"01000101", 
"10001100", 
"10011001", 
"01111010", 
"10010010", 
"10001010", 
"01100001", 
"10001000", 
"01010100", 
"01000011", 
"01011101", 
"01010010", 
"01111010", 
"10010101", 
"10101110", 
"10001101", 
"01100101", 
"10000011", 
"10000001", 
"01101110", 
"01111010", 
"10100001", 
"10000010", 
"01100110", 
"01110111", 
"01010010", 
"10000010", 
"01110110", 
"10001011", 
"10001101", 
"10011010", 
"10100101", 
"01100011", 
"10010001", 
"01111101", 
"01101000", 
"10110001", 
"01110011", 
"01111101", 
"01111111", 
"10000000", 
"10100011", 
"01000111", 
"01101100", 
"10111001", 
"10010011", 
"10000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_45: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_45(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
