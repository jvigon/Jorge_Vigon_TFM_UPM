use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_1_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_1_LAYER;

architecture Behavioral of ROM_FC_84_1_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_1: ROM_ARRAY_PESOS_FC_84 := (
"01111111", 
"01111011", 
"10000110", 
"10001001", 
"01110110", 
"10001000", 
"10000101", 
"01000111", 
"01101001", 
"10011111", 
"01101110", 
"10100000", 
"01101111", 
"01101101", 
"01100010", 
"01110011", 
"01101110", 
"10100010", 
"10010001", 
"10101101", 
"01110010", 
"01001011", 
"01110101", 
"01111001", 
"10001011", 
"10010000", 
"01110101", 
"10000111", 
"10010001", 
"01010100", 
"01110110", 
"01111111", 
"10001001", 
"01101010", 
"10001000", 
"10101100", 
"01110010", 
"10000001", 
"01111101", 
"01101100", 
"10001110", 
"01111101", 
"01011011", 
"01011001", 
"10001111", 
"01010111", 
"01110011", 
"10001011", 
"01110001", 
"10000010", 
"01110011", 
"10001011", 
"10010011", 
"01100111", 
"01000010", 
"01100011", 
"10010000", 
"01101100", 
"10001000", 
"01111000", 
"01110110", 
"01011010", 
"01011110", 
"01110001", 
"10001011", 
"10001000", 
"10010011", 
"10010000", 
"10001001", 
"01100101", 
"01111010", 
"01011010", 
"10000010", 
"10101010", 
"10001001", 
"10000011", 
"01100011", 
"10011100", 
"01101111", 
"01011011", 
"01100101", 
"10100011", 
"10001110", 
"01011100", 
"10010101", 
"10001101", 
"01101110", 
"10001000", 
"01111110", 
"01111000", 
"10011101", 
"01100111", 
"01101110", 
"10001111", 
"01111011", 
"10000011", 
"01110101", 
"10001010", 
"10000011", 
"10001010", 
"10001010", 
"01110101", 
"10110101", 
"01001110", 
"10010100", 
"01111100", 
"10010000", 
"10001101", 
"01110001", 
"01011011", 
"10010101", 
"10000100", 
"10010101", 
"10000010", 
"10010000", 
"10010111", 
"10001101", 
"01101011", 
"10010110", 
"01101100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_1 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_1(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
