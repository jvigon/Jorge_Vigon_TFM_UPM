use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_14_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_14_LAYER;

architecture Behavioral of ROM_FC_84_14_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_14: ROM_ARRAY_PESOS_FC_84 := (
"01110011", 
"01101110", 
"10000011", 
"10001011", 
"10000011", 
"01101010", 
"01111100", 
"10010011", 
"01000111", 
"01101101", 
"10001101", 
"10010111", 
"01101011", 
"10001000", 
"10011001", 
"10101011", 
"01010000", 
"10010100", 
"01101000", 
"00111100", 
"10100010", 
"01000001", 
"10010100", 
"01011011", 
"01111010", 
"10000110", 
"01101101", 
"10000000", 
"01110110", 
"10100010", 
"01111011", 
"01101001", 
"01111111", 
"10101101", 
"01011110", 
"10010111", 
"01100100", 
"01101101", 
"10011110", 
"10000101", 
"10010110", 
"01111011", 
"01000010", 
"10001010", 
"10101100", 
"01110011", 
"01110111", 
"01110110", 
"01100100", 
"01111011", 
"01111011", 
"11010001", 
"10000110", 
"01110111", 
"01111111", 
"10000000", 
"10010101", 
"10000010", 
"01111010", 
"10001010", 
"01101001", 
"01011110", 
"10100010", 
"01010010", 
"01010000", 
"01100001", 
"01111010", 
"01110011", 
"10011101", 
"10010001", 
"01010001", 
"01000010", 
"01111101", 
"01100010", 
"01101011", 
"10001110", 
"01111100", 
"01100011", 
"01110100", 
"01010011", 
"01111101", 
"10010101", 
"01100010", 
"01000100", 
"01011001", 
"01111001", 
"10001100", 
"01001110", 
"01110000", 
"01100100", 
"01001110", 
"01111111", 
"10001110", 
"01100000", 
"01101111", 
"10100000", 
"01100010", 
"10001100", 
"01011011", 
"01111010", 
"10000110", 
"01110110", 
"01100000", 
"01100111", 
"01001110", 
"10011101", 
"01110111", 
"01101110", 
"01111000", 
"10010011", 
"10100101", 
"10000010", 
"01110110", 
"01010100", 
"01111100", 
"01111101", 
"10010011", 
"01010110", 
"10000010", 
"10011011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_14 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_14(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
