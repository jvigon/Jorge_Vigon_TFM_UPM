use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_32_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_32_LAYER;

architecture Behavioral of ROM_FC_84_32_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_32: ROM_ARRAY_PESOS_FC_84 := (
"01111010", 
"01100000", 
"01110101", 
"10011101", 
"01110100", 
"01100001", 
"10001011", 
"01101011", 
"10011001", 
"10000101", 
"10011100", 
"01011110", 
"01011100", 
"01101011", 
"10110010", 
"10000011", 
"01111110", 
"10010011", 
"01100100", 
"10000111", 
"10010001", 
"10001011", 
"01101110", 
"01111001", 
"10011000", 
"01110010", 
"01011001", 
"01101101", 
"10000100", 
"10001001", 
"10001110", 
"01111011", 
"10001101", 
"01100001", 
"01110111", 
"01011010", 
"01111110", 
"10010011", 
"10100010", 
"10010110", 
"01011101", 
"01111000", 
"01101010", 
"01100100", 
"01011011", 
"01011010", 
"01011111", 
"10010100", 
"01010000", 
"10010000", 
"01100001", 
"01111110", 
"10011000", 
"10000000", 
"01100100", 
"10100110", 
"01101100", 
"01100110", 
"01111000", 
"01101111", 
"01100001", 
"01010000", 
"10000100", 
"01111101", 
"01111110", 
"01011101", 
"01111000", 
"01101110", 
"01100101", 
"10010111", 
"01010001", 
"01101110", 
"01001101", 
"01011101", 
"01110001", 
"10010000", 
"01011111", 
"01111001", 
"01111101", 
"01101011", 
"10001100", 
"01011110", 
"01001110", 
"01101110", 
"10000001", 
"01110001", 
"01101110", 
"01011110", 
"01110001", 
"10000101", 
"01110111", 
"10011111", 
"10001000", 
"01110010", 
"01001010", 
"01100011", 
"10001011", 
"10010100", 
"01111111", 
"10000011", 
"10010001", 
"10010100", 
"01010011", 
"01100111", 
"10001001", 
"01101001", 
"01101101", 
"01110010", 
"01010101", 
"10001110", 
"10001010", 
"10001000", 
"10010010", 
"01111010", 
"01101011", 
"10001100", 
"01101000", 
"01111100", 
"01111001", 
"01011001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_32 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_32(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
