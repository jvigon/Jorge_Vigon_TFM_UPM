use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_31_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_31_LAYER;

architecture Behavioral of ROM_FC_84_31_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_31: ROM_ARRAY_PESOS_FC_84 := (
"01110100", 
"01111101", 
"10010011", 
"10001011", 
"10010100", 
"10000110", 
"10010111", 
"01110110", 
"10110011", 
"10011000", 
"10000000", 
"10000101", 
"01100110", 
"01110000", 
"10001111", 
"01100101", 
"01111100", 
"01110011", 
"01101010", 
"01101000", 
"10101101", 
"10010011", 
"10000010", 
"01111001", 
"01101100", 
"01111001", 
"10011010", 
"10000100", 
"01011011", 
"10001011", 
"01100110", 
"01100000", 
"01100111", 
"01100010", 
"00101011", 
"10100110", 
"01011110", 
"10000101", 
"01110010", 
"01100100", 
"10010000", 
"10001010", 
"01101011", 
"01100100", 
"01101001", 
"01111110", 
"10010011", 
"01000011", 
"01111011", 
"10000100", 
"10001001", 
"01110110", 
"10100000", 
"10001110", 
"01111111", 
"01111010", 
"10010010", 
"01111001", 
"10101000", 
"01110011", 
"10001100", 
"10011000", 
"01110110", 
"10011001", 
"01001011", 
"10111011", 
"01000101", 
"01111010", 
"10001111", 
"01010010", 
"01110000", 
"10100010", 
"10100111", 
"01111101", 
"10011011", 
"10001000", 
"10001011", 
"10000010", 
"10011110", 
"01000000", 
"01111011", 
"10010000", 
"01110100", 
"01000101", 
"10000010", 
"01100010", 
"01010010", 
"01101111", 
"01111010", 
"01001110", 
"10000101", 
"10010000", 
"01110001", 
"01001001", 
"10001010", 
"10010001", 
"01011110", 
"01111101", 
"10110011", 
"01100101", 
"10011000", 
"01110110", 
"01101100", 
"01010010", 
"00101111", 
"01110000", 
"01100110", 
"01111010", 
"00110101", 
"01100011", 
"01000101", 
"10010111", 
"01100010", 
"01001101", 
"01101100", 
"01011100", 
"10001001", 
"10001000", 
"10010011", 
"01100000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_31 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_31(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
