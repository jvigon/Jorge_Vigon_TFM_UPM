use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_41_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_41_LAYER;

architecture Behavioral of ROM_FC_84_41_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_41: ROM_ARRAY_PESOS_FC_84 := (
"01101100", 
"01111101", 
"10101100", 
"10010110", 
"01100110", 
"01101111", 
"10000111", 
"10000010", 
"01101001", 
"10000111", 
"10011101", 
"01011100", 
"10001101", 
"10100111", 
"11000101", 
"10000101", 
"10100001", 
"10100001", 
"10010000", 
"10001001", 
"01110010", 
"10011110", 
"10010101", 
"01101010", 
"01111101", 
"10101110", 
"01110110", 
"10010011", 
"01100110", 
"10100010", 
"01101110", 
"01011101", 
"10010101", 
"10001110", 
"01001111", 
"01100101", 
"10001011", 
"01010101", 
"10011010", 
"01101010", 
"01000111", 
"01110110", 
"01011010", 
"01010111", 
"10010111", 
"10100001", 
"01010110", 
"10001001", 
"00111011", 
"01101011", 
"01101101", 
"01111101", 
"10000010", 
"01101001", 
"10011101", 
"01011110", 
"01100011", 
"01100000", 
"01110101", 
"10010001", 
"10011000", 
"10010011", 
"01111011", 
"01010111", 
"01110110", 
"01111110", 
"10001110", 
"01110111", 
"10000001", 
"10001101", 
"01100011", 
"01000101", 
"01110101", 
"01011111", 
"01011111", 
"10010111", 
"10011001", 
"10000011", 
"10011010", 
"10000110", 
"01101010", 
"01110010", 
"10001111", 
"01111101", 
"01000111", 
"01011001", 
"01111111", 
"01001010", 
"10010110", 
"01010001", 
"01111110", 
"10001000", 
"10011101", 
"01100001", 
"10000001", 
"01111100", 
"01111101", 
"10011100", 
"10000011", 
"10011011", 
"10000011", 
"10010100", 
"01100110", 
"01100011", 
"01010110", 
"01110101", 
"10000111", 
"01111010", 
"10000000", 
"10101100", 
"01111100", 
"10000100", 
"10001001", 
"10100010", 
"01110000", 
"10010010", 
"01111111", 
"01111000", 
"10001100", 
"01010110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_41: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_41(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
