use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_44_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_44_LAYER;

architecture Behavioral of ROM_FC_84_44_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_44: ROM_ARRAY_PESOS_FC_84 := (
"01000100", 
"01100000", 
"01101010", 
"10010011", 
"10000101", 
"10110010", 
"01101001", 
"01110010", 
"10001101", 
"10110010", 
"10100100", 
"10010011", 
"10000110", 
"01110111", 
"01110100", 
"10010001", 
"10010101", 
"01100111", 
"01110000", 
"01100111", 
"01111111", 
"00111100", 
"10100011", 
"10100000", 
"01111111", 
"10011101", 
"01110011", 
"10001111", 
"01100111", 
"01101011", 
"01111110", 
"10000010", 
"10001011", 
"10010010", 
"01010011", 
"01110100", 
"01100111", 
"10000100", 
"10011010", 
"10100101", 
"01110101", 
"00111001", 
"01100001", 
"10100010", 
"10100101", 
"00111100", 
"10100101", 
"01111010", 
"10000000", 
"10001101", 
"10101110", 
"10000101", 
"10001001", 
"10000111", 
"10011001", 
"10010010", 
"10000101", 
"01101110", 
"10001001", 
"01001110", 
"01101000", 
"10010110", 
"10001100", 
"10001100", 
"01111100", 
"10001001", 
"10101000", 
"10010001", 
"10000111", 
"10000010", 
"01101111", 
"01100000", 
"01100010", 
"01011111", 
"10000010", 
"01110010", 
"10011000", 
"01111010", 
"10000011", 
"10000000", 
"10000101", 
"10010100", 
"10010000", 
"01101000", 
"10000011", 
"10011111", 
"10010011", 
"01011010", 
"01101100", 
"10000110", 
"01110100", 
"01010010", 
"01111001", 
"01111101", 
"01100110", 
"01111000", 
"01101111", 
"01100100", 
"10001100", 
"10010100", 
"01111001", 
"10001000", 
"10000101", 
"10000010", 
"01100000", 
"10001101", 
"01110111", 
"10011010", 
"01001011", 
"01001111", 
"10000000", 
"10001000", 
"01110001", 
"01010110", 
"10001001", 
"10010101", 
"10101111", 
"01101000", 
"10001001", 
"01101111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_44: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_44(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
