use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_61_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_61_LAYER;

architecture Behavioral of ROM_FC_84_61_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_61: ROM_ARRAY_PESOS_FC_84 := (
"10001010", 
"01101111", 
"01100011", 
"10010111", 
"01101110", 
"01101111", 
"10010000", 
"01100110", 
"00111110", 
"01110000", 
"01011100", 
"01110010", 
"10010010", 
"01101101", 
"10001010", 
"01110100", 
"01110001", 
"10011001", 
"10000101", 
"10001100", 
"01111010", 
"01101011", 
"10001101", 
"01100010", 
"10011111", 
"10011110", 
"01101101", 
"01011101", 
"10001010", 
"01100001", 
"10010010", 
"01000110", 
"10100110", 
"01110010", 
"01100110", 
"01100101", 
"10010011", 
"01110100", 
"01110111", 
"01111000", 
"10001010", 
"01011101", 
"01111010", 
"10011010", 
"01111010", 
"01100101", 
"01110000", 
"01101011", 
"01101101", 
"10011101", 
"10000111", 
"10011101", 
"01101100", 
"10000011", 
"01100101", 
"10000101", 
"01111000", 
"10011000", 
"10000010", 
"10001011", 
"01110001", 
"01100011", 
"10001011", 
"10010010", 
"10000101", 
"01011111", 
"10100110", 
"10000011", 
"01100111", 
"01110011", 
"01111011", 
"01110110", 
"01001011", 
"10000110", 
"10011111", 
"01101001", 
"01100000", 
"10001101", 
"01110000", 
"01101011", 
"10001001", 
"01111010", 
"10010010", 
"01011111", 
"01011011", 
"10000000", 
"10011001", 
"01111110", 
"10011000", 
"01100001", 
"10110110", 
"10010100", 
"01111100", 
"01100110", 
"01010000", 
"10001101", 
"01011101", 
"01110000", 
"10001001", 
"01111101", 
"01011100", 
"10010001", 
"10011101", 
"01111110", 
"10001000", 
"10011001", 
"01110001", 
"10100011", 
"10011010", 
"01110001", 
"01011101", 
"01011101", 
"01111100", 
"00111001", 
"01101011", 
"10010011", 
"01110011", 
"01111001", 
"10000101", 
"01110111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_61 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_61(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
