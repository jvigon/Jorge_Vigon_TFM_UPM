use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_4_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_4_LAYER;

architecture Behavioral of ROM_FC_84_4_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_4: ROM_ARRAY_PESOS_FC_84 := (
"01110111", 
"10010011", 
"01100101", 
"10010000", 
"01011000", 
"10011011", 
"01101001", 
"01011100", 
"01101001", 
"10100100", 
"10001010", 
"00111101", 
"00110111", 
"01111110", 
"00111001", 
"01011111", 
"10100000", 
"10001100", 
"10000111", 
"11001010", 
"01111000", 
"01111100", 
"01011010", 
"01110110", 
"10011000", 
"00110110", 
"01001111", 
"10010010", 
"01111100", 
"10001101", 
"10011001", 
"10000010", 
"01110101", 
"01011100", 
"01111100", 
"01000111", 
"01111011", 
"01100100", 
"01111110", 
"01111010", 
"10001100", 
"01110111", 
"01110011", 
"10000000", 
"01001001", 
"01011100", 
"01000101", 
"10001010", 
"01011010", 
"01110010", 
"01111010", 
"10010010", 
"01101100", 
"01011001", 
"01110001", 
"10111100", 
"10001110", 
"10001010", 
"01111001", 
"10001101", 
"01010100", 
"01100111", 
"01110000", 
"01011001", 
"11001010", 
"00111011", 
"10011100", 
"10011110", 
"01111001", 
"01100110", 
"01111001", 
"01010111", 
"10001010", 
"10101011", 
"10000101", 
"10001101", 
"01011100", 
"01101110", 
"00111010", 
"01011010", 
"01100101", 
"00111000", 
"01100110", 
"10010100", 
"01000111", 
"10000011", 
"01100101", 
"10000100", 
"10001111", 
"01110001", 
"00111101", 
"10111111", 
"01110111", 
"01110011", 
"01111000", 
"01110010", 
"10011010", 
"01101011", 
"01001101", 
"10000100", 
"01100111", 
"01100011", 
"01110001", 
"01111010", 
"01111011", 
"10001100", 
"10000111", 
"01111011", 
"10100100", 
"01111101", 
"10101100", 
"10001000", 
"10000110", 
"10011001", 
"01101110", 
"10000100", 
"01111000", 
"10000111", 
"01101111", 
"10110011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_4 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_4(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
