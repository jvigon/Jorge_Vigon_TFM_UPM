use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_68_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_68_LAYER;

architecture Behavioral of ROM_FC_84_68_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_68: ROM_ARRAY_PESOS_FC_84 := (
"10001001", 
"01001111", 
"10001110", 
"10011101", 
"10000101", 
"10001100", 
"01111000", 
"10001010", 
"01100010", 
"01100010", 
"01110010", 
"10000000", 
"01110111", 
"01111111", 
"01100011", 
"10010011", 
"10001010", 
"01011011", 
"01111100", 
"01101010", 
"10001000", 
"01100011", 
"10010011", 
"01110110", 
"01110001", 
"10000011", 
"01001101", 
"10000111", 
"10011110", 
"01101010", 
"10101111", 
"10001000", 
"00110100", 
"01000100", 
"10101111", 
"01111001", 
"01111101", 
"01111100", 
"10011000", 
"01100010", 
"01001001", 
"10001010", 
"10010010", 
"01100010", 
"01101111", 
"01100000", 
"10001110", 
"10000000", 
"10100011", 
"01101111", 
"01011011", 
"01110010", 
"10000101", 
"10100000", 
"00111100", 
"10000000", 
"01100011", 
"01110101", 
"01100111", 
"10011001", 
"10001111", 
"01010011", 
"10000110", 
"01001101", 
"10100101", 
"00101111", 
"10000100", 
"10011111", 
"10000011", 
"01101000", 
"01110100", 
"01100111", 
"10000111", 
"01100101", 
"10011110", 
"01110100", 
"01101001", 
"10000100", 
"10000101", 
"10010000", 
"10010101", 
"10011110", 
"01000010", 
"01111100", 
"10000111", 
"01011110", 
"10011011", 
"01110000", 
"10000101", 
"10101001", 
"01101111", 
"10010110", 
"01001100", 
"10000001", 
"01101111", 
"01110011", 
"01110010", 
"10011100", 
"10000100", 
"01100101", 
"10000110", 
"10010111", 
"01101011", 
"01101010", 
"10100101", 
"10011011", 
"01101100", 
"01110110", 
"01110110", 
"01000010", 
"01111011", 
"01111100", 
"01110011", 
"10011011", 
"01101110", 
"10001010", 
"10010101", 
"10011011", 
"01110000", 
"01100010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_68: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_68(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
