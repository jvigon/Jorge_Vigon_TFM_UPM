use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_57_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_57_LAYER;

architecture Behavioral of ROM_FC_84_57_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_57: ROM_ARRAY_PESOS_FC_84 := (
"10001111", 
"01111111", 
"01010000", 
"10000111", 
"10001110", 
"01111101", 
"10010000", 
"00111001", 
"01100001", 
"01101111", 
"10010110", 
"01001100", 
"01001010", 
"10100001", 
"01011110", 
"10010110", 
"01101010", 
"10101000", 
"01101001", 
"01110101", 
"10100101", 
"10001011", 
"10010100", 
"01001110", 
"01111111", 
"01100111", 
"01001000", 
"01111000", 
"10001001", 
"01100000", 
"01101101", 
"01010100", 
"01110011", 
"10100001", 
"01001101", 
"01001101", 
"01111011", 
"01011000", 
"01111110", 
"10010011", 
"10000100", 
"01101001", 
"10100110", 
"10000111", 
"01101011", 
"01101110", 
"01100001", 
"10011011", 
"01011110", 
"10011001", 
"01101011", 
"10001111", 
"01111111", 
"01110011", 
"01001010", 
"10001100", 
"10001001", 
"01101010", 
"01011010", 
"01101100", 
"10001110", 
"10000110", 
"10011010", 
"01001111", 
"10000000", 
"01101011", 
"01111100", 
"10001111", 
"01111100", 
"10010011", 
"01101000", 
"10000011", 
"10001111", 
"01101111", 
"01110000", 
"10010000", 
"01001000", 
"01101110", 
"01110100", 
"01011001", 
"01011001", 
"01011110", 
"01010010", 
"01010111", 
"01101100", 
"10010010", 
"01111100", 
"01011001", 
"10010001", 
"01000110", 
"01011100", 
"10011111", 
"10010010", 
"10000110", 
"00111111", 
"01110110", 
"01110100", 
"10100101", 
"01111111", 
"10001011", 
"10010100", 
"01100110", 
"01111110", 
"01101010", 
"10110110", 
"01101110", 
"10001101", 
"10010000", 
"01111001", 
"10001111", 
"01111101", 
"01111101", 
"10011000", 
"10010010", 
"10011001", 
"10100100", 
"01100100", 
"10101100", 
"01101010", 
"10010101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_57 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_57(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
