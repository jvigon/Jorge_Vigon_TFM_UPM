use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_13_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_13_LAYER;

architecture Behavioral of ROM_FC_120_13_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_13: ROM_ARRAY_PESOS_FC_120 := (
"10011001", 
"01000011", 
"01110010", 
"10011001", 
"10001010", 
"10100010", 
"01010100", 
"01101110", 
"01100100", 
"01110011", 
"10101010", 
"01101110", 
"01111101", 
"10110111", 
"01111010", 
"10010000", 
"10001011", 
"00110101", 
"01010011", 
"01101011", 
"01111000", 
"01100001", 
"01101111", 
"10100010", 
"01110111", 
"01011011", 
"01000100", 
"01111010", 
"01011011", 
"10000100", 
"10000101", 
"01111110", 
"01110111", 
"01011001", 
"01100011", 
"01011100", 
"10010000", 
"01101011", 
"10011001", 
"01111110", 
"01101110", 
"01110100", 
"01110111", 
"10000010", 
"10101011", 
"01110100", 
"10011000", 
"10010011", 
"10001000", 
"01111101", 
"10000000", 
"01000011", 
"01111100", 
"10000001", 
"10001101", 
"10000001", 
"01110000", 
"01111101", 
"01010110", 
"10100100", 
"10011011", 
"01010100", 
"01110110", 
"10110101", 
"01011101", 
"01101000", 
"10110011", 
"10011100", 
"10000100", 
"10101010", 
"00111101", 
"01101110", 
"01111000", 
"01111101", 
"10111001", 
"01011111", 
"01111101", 
"11000111", 
"10001100", 
"01110111", 
"01000011", 
"01100111", 
"10000010", 
"10101000", 
"01110110", 
"01101010", 
"10000111", 
"10000011", 
"01101110", 
"01111001", 
"01110110", 
"01010011", 
"01101100", 
"10110110", 
"10010111", 
"10001010", 
"01011101", 
"01011010", 
"01100111", 
"01110110", 
"10100101", 
"01111100", 
"01111011", 
"01011101", 
"01101011", 
"01111010", 
"01111111", 
"01111001", 
"01110010", 
"01101000", 
"10011000", 
"01110001", 
"01101011", 
"01100000", 
"10100001", 
"10010110", 
"01101101", 
"01110011", 
"01101011", 
"01101100", 
"01110001", 
"01101110", 
"10001000", 
"01011100", 
"01011010", 
"10000010", 
"10001100", 
"10111001", 
"01010101", 
"01100001", 
"10000111", 
"01101101", 
"01100010", 
"10001110", 
"01011111", 
"10001011", 
"10010000", 
"01101101", 
"10101010", 
"01100101", 
"01100011", 
"10011010", 
"10000001", 
"10001010", 
"01110011", 
"01111010", 
"10000000", 
"01101100", 
"01111111", 
"01110001", 
"01011000", 
"01010010", 
"01101101", 
"01001101", 
"01101101", 
"01101101", 
"01111101", 
"10110010", 
"01110000", 
"01111100", 
"10010010", 
"01010110", 
"01111100", 
"10001001", 
"01111100", 
"01111110", 
"01100101", 
"01111000", 
"10000111", 
"01111100", 
"10000000", 
"01010010", 
"01110101", 
"01100101", 
"10000011", 
"01110011", 
"01100010", 
"01000101", 
"10000101", 
"11000100", 
"01101111", 
"01101101", 
"01010011", 
"01100001", 
"01110011", 
"10100100", 
"01111011", 
"01000010", 
"01110010", 
"01000111", 
"01111011", 
"01110100", 
"01101001", 
"10100110", 
"01101000", 
"01010100", 
"01111001", 
"01101110", 
"01111100", 
"01101101", 
"10010000", 
"01110011", 
"10000010", 
"01011011", 
"01011111", 
"10001101", 
"01111111", 
"01110110", 
"01100010", 
"10000100", 
"01101100", 
"10000001", 
"10001111", 
"01101010", 
"01110100", 
"01100001", 
"10010010", 
"10000101", 
"01101010", 
"01111001", 
"01011100", 
"10010011", 
"01101011", 
"10001110", 
"01100110", 
"01110011", 
"10001101", 
"10000001", 
"10000100", 
"01110101", 
"01101000", 
"10000110", 
"10001010", 
"10010000", 
"10001111", 
"01011100", 
"10001110", 
"10010011", 
"10001001", 
"01111010", 
"01101001", 
"01100101", 
"01111010", 
"01000111", 
"01110100", 
"01000111", 
"01111010", 
"01101000", 
"10010001", 
"10001011", 
"01110011", 
"01010001", 
"01001000", 
"10000110", 
"01100100", 
"01101101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_13: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_13(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
