use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_65_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_65_LAYER;

architecture Behavioral of ROM_FC_120_65_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_65: ROM_ARRAY_PESOS_FC_120 := (
"01111010", 
"01001001", 
"10011001", 
"10111011", 
"01011111", 
"10000011", 
"10101011", 
"01101111", 
"10000001", 
"10010010", 
"10011000", 
"10000000", 
"10100110", 
"10010011", 
"01101110", 
"10001011", 
"10011000", 
"10001100", 
"10011110", 
"10100011", 
"01101111", 
"01011110", 
"01010011", 
"10000001", 
"10000001", 
"10001000", 
"10000000", 
"10011111", 
"10100101", 
"01010011", 
"01110100", 
"10000011", 
"10010100", 
"01110101", 
"01100101", 
"10001100", 
"01100111", 
"01111010", 
"01000110", 
"01110011", 
"10001000", 
"11000010", 
"01100111", 
"10010000", 
"10011100", 
"01111111", 
"01110101", 
"01101111", 
"10100100", 
"10001010", 
"01010101", 
"01011011", 
"01111000", 
"01101000", 
"01111011", 
"01011110", 
"01111001", 
"10111010", 
"01111110", 
"10100110", 
"10100111", 
"01001011", 
"01111011", 
"10001100", 
"01110111", 
"10001101", 
"10000100", 
"10000010", 
"10000110", 
"01110011", 
"10001010", 
"01000011", 
"10001010", 
"10001111", 
"01011111", 
"01111011", 
"10001101", 
"10000101", 
"10000011", 
"01111001", 
"01110101", 
"10000101", 
"10001111", 
"10100011", 
"10100100", 
"01011101", 
"10011011", 
"01011110", 
"01101111", 
"10001100", 
"10000001", 
"10001110", 
"10010001", 
"10010111", 
"10001100", 
"01101001", 
"10010111", 
"01111101", 
"10010100", 
"10110101", 
"10001011", 
"10000000", 
"01011100", 
"01100000", 
"10001100", 
"10010001", 
"00111001", 
"10010010", 
"10001010", 
"01110111", 
"10000100", 
"01110110", 
"10011001", 
"01110100", 
"10001011", 
"01110100", 
"01110111", 
"01110010", 
"01000001", 
"01111101", 
"01101011", 
"10100000", 
"01111011", 
"10100011", 
"10000011", 
"01110101", 
"01110011", 
"01111001", 
"01110001", 
"10110000", 
"00101101", 
"01101000", 
"01111000", 
"01110110", 
"10010101", 
"01111010", 
"10000101", 
"01110100", 
"01011110", 
"10101101", 
"01101110", 
"01101010", 
"01111011", 
"10010010", 
"01010100", 
"01111011", 
"01101100", 
"10001100", 
"01100110", 
"10011110", 
"10101110", 
"10001100", 
"10000011", 
"01110000", 
"01111110", 
"01011111", 
"01111100", 
"01110110", 
"10000101", 
"01100110", 
"10010101", 
"01110011", 
"01110111", 
"01111111", 
"10000011", 
"01100010", 
"01010110", 
"01110111", 
"10000111", 
"10010011", 
"01110111", 
"10000000", 
"01111010", 
"01011000", 
"01101110", 
"10000100", 
"10011001", 
"10100011", 
"10010000", 
"10010111", 
"01111111", 
"01001010", 
"01010110", 
"01111000", 
"10000111", 
"01101001", 
"01110001", 
"10110011", 
"00011101", 
"10100111", 
"10000001", 
"01100110", 
"01101110", 
"10111011", 
"01110010", 
"01110101", 
"10001111", 
"01101101", 
"10101011", 
"01110010", 
"01110000", 
"00110000", 
"01011101", 
"11010100", 
"10000111", 
"01001110", 
"10010011", 
"01110011", 
"01101101", 
"10100010", 
"10001100", 
"01101011", 
"10001100", 
"10001011", 
"10000100", 
"10000101", 
"10001010", 
"01100011", 
"10111011", 
"01000011", 
"01101001", 
"01010000", 
"10010000", 
"10001010", 
"10011100", 
"10100111", 
"01101011", 
"10000011", 
"10011010", 
"10100011", 
"01101010", 
"10011000", 
"01110011", 
"01110110", 
"10111010", 
"01001100", 
"01011000", 
"01100010", 
"01111001", 
"10001100", 
"01111111", 
"10110100", 
"01100111", 
"01001110", 
"10001111", 
"10001111", 
"10010001", 
"10010001", 
"10001000", 
"01010000", 
"01100101", 
"10000001", 
"01111011", 
"01101010", 
"10010000", 
"01110101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_65: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_65(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
