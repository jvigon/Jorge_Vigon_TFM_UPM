use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_2_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_2_LAYER;

architecture Behavioral of ROM_FC_120_2_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_2: ROM_ARRAY_PESOS_FC_120 := (
"01111100", 
"10001101", 
"00101101", 
"01001001", 
"10100100", 
"10101001", 
"10000111", 
"01110011", 
"01111100", 
"00101001", 
"01001000", 
"01010010", 
"01110000", 
"01111110", 
"01111111", 
"01100010", 
"01110001", 
"01111101", 
"01100001", 
"01110100", 
"01100111", 
"10100011", 
"10001010", 
"01110111", 
"10000000", 
"00111000", 
"01011000", 
"00110000", 
"01010010", 
"10011110", 
"01111000", 
"01111100", 
"10010101", 
"01001101", 
"01011001", 
"01111101", 
"10011000", 
"10010011", 
"10111110", 
"10010100", 
"10000101", 
"01110001", 
"10100000", 
"01011010", 
"01011100", 
"10010000", 
"10000111", 
"01101000", 
"10110011", 
"01110111", 
"10001010", 
"01111001", 
"10001100", 
"10010000", 
"10100111", 
"01110000", 
"10001010", 
"10010000", 
"01111000", 
"10000011", 
"01101100", 
"10000000", 
"10010100", 
"01110111", 
"01110010", 
"10010101", 
"10011010", 
"10011111", 
"01100011", 
"10000100", 
"01101111", 
"01101000", 
"01101111", 
"01010010", 
"01100110", 
"01011011", 
"10010111", 
"10010001", 
"01111000", 
"01111010", 
"01100100", 
"01111001", 
"10011010", 
"10001010", 
"01111001", 
"10001010", 
"01110100", 
"10010010", 
"01010101", 
"01000001", 
"01100100", 
"00101000", 
"01110011", 
"01000110", 
"10001001", 
"01101011", 
"10011111", 
"01011011", 
"01110001", 
"10000000", 
"10000000", 
"10010000", 
"01101110", 
"10000011", 
"10100110", 
"10010110", 
"10011010", 
"01101001", 
"01010111", 
"10010101", 
"01110001", 
"10000100", 
"10001100", 
"01000000", 
"01101100", 
"10000110", 
"01100011", 
"01110101", 
"01111001", 
"10010101", 
"01101100", 
"01111101", 
"10010100", 
"01100111", 
"10100010", 
"01100100", 
"10001000", 
"10001000", 
"10010100", 
"01111100", 
"00000100", 
"01110010", 
"01111000", 
"10000110", 
"10000110", 
"10001110", 
"10000111", 
"10110110", 
"01010110", 
"10000000", 
"01010100", 
"00111000", 
"10000001", 
"01100000", 
"10011011", 
"01111010", 
"01011110", 
"01001010", 
"01111011", 
"10010011", 
"01110111", 
"10001001", 
"01110110", 
"01110000", 
"01010001", 
"01010001", 
"01011001", 
"01010111", 
"10010001", 
"01100011", 
"10101010", 
"01100010", 
"01000001", 
"10000111", 
"01111100", 
"10010000", 
"01101001", 
"10100000", 
"10010011", 
"01101111", 
"10010000", 
"01101011", 
"01011100", 
"10101000", 
"10010110", 
"01101110", 
"01101001", 
"01101100", 
"01111000", 
"01100000", 
"10000101", 
"01101110", 
"01100000", 
"10000101", 
"01101110", 
"01001101", 
"01110001", 
"01111110", 
"01100100", 
"10011100", 
"10000111", 
"01110111", 
"10101111", 
"01011110", 
"01110111", 
"10001001", 
"01110010", 
"10011100", 
"01111011", 
"10100001", 
"01111111", 
"01111010", 
"10000100", 
"10110011", 
"01111000", 
"01000011", 
"10000001", 
"10001010", 
"10001011", 
"10010000", 
"01110001", 
"01100100", 
"01110110", 
"10101100", 
"00111000", 
"10000100", 
"01101101", 
"01011000", 
"10001001", 
"01111110", 
"01101110", 
"01101101", 
"10001110", 
"10000000", 
"01111111", 
"10000000", 
"10011110", 
"10010001", 
"01111001", 
"01110101", 
"01111101", 
"10101010", 
"01011000", 
"01011101", 
"01101111", 
"01001111", 
"01111001", 
"10001010", 
"01111100", 
"10000110", 
"01110011", 
"10101011", 
"10001110", 
"10010101", 
"10001110", 
"10010100", 
"10000010", 
"01111001", 
"10000111", 
"01101001", 
"10000100", 
"01010111", 
"10101011", 
"10001001", 
"10010000", 
"10011010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_2 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_2(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
