use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_11_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_11_LAYER;

architecture Behavioral of ROM_FC_84_11_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_11: ROM_ARRAY_PESOS_FC_84 := (
"10000110", 
"01110011", 
"10001000", 
"01111010", 
"01111010", 
"10011011", 
"01111011", 
"01111100", 
"10011000", 
"10001010", 
"10011010", 
"10001001", 
"01001101", 
"10011000", 
"01001001", 
"01011100", 
"10010001", 
"10011110", 
"01101000", 
"01101010", 
"01100111", 
"01101010", 
"10000010", 
"01010111", 
"01011111", 
"01111001", 
"01110011", 
"01110011", 
"01001011", 
"01110101", 
"01111011", 
"01011110", 
"10100100", 
"10011011", 
"01100111", 
"01001101", 
"01101010", 
"01110110", 
"00111001", 
"01111000", 
"01111111", 
"01011101", 
"01110011", 
"10011001", 
"01100001", 
"01111000", 
"10001110", 
"10010110", 
"01100011", 
"01110001", 
"01110100", 
"01111101", 
"10000001", 
"10010010", 
"10010010", 
"01011000", 
"10010010", 
"10000000", 
"01100100", 
"01100111", 
"01011110", 
"10000101", 
"01111010", 
"10000001", 
"10001000", 
"10010001", 
"10011100", 
"01101001", 
"10010000", 
"10110001", 
"01011101", 
"01110101", 
"01101010", 
"01101011", 
"10001101", 
"10010011", 
"01100100", 
"10001011", 
"01101011", 
"01010000", 
"01101110", 
"10000001", 
"01110101", 
"01010010", 
"01011000", 
"01011110", 
"00110011", 
"01100111", 
"01101011", 
"01111110", 
"01101001", 
"01101000", 
"01111100", 
"01010110", 
"01011101", 
"01111010", 
"01010100", 
"01101001", 
"01100001", 
"01100100", 
"10001010", 
"01111101", 
"01101110", 
"00111110", 
"01111010", 
"01101100", 
"01110001", 
"01101111", 
"01011000", 
"01111110", 
"01101011", 
"01111100", 
"10001000", 
"01101001", 
"10010001", 
"10100001", 
"01110111", 
"01010101", 
"01110010", 
"01011000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_11 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_11(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
