use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_0_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_0_LAYER;

architecture Behavioral of ROM_FC_84_0_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_0: ROM_ARRAY_PESOS_FC_84 := (
"10100011", 
"10100100", 
"01011000", 
"01110010", 
"01100000", 
"01100110", 
"10010010", 
"01001101", 
"10100010", 
"11000100", 
"01110000", 
"01111011", 
"00111011", 
"01101101", 
"01101001", 
"01101111", 
"01110100", 
"01111010", 
"01100000", 
"01110010", 
"01101001", 
"01011111", 
"10000100", 
"10000110", 
"01110111", 
"10001110", 
"10010110", 
"10011110", 
"10100100", 
"01110111", 
"10011001", 
"10010101", 
"10100000", 
"10011110", 
"01011010", 
"10000110", 
"01111100", 
"01111001", 
"01101110", 
"01110001", 
"01001110", 
"01111010", 
"01000001", 
"00011011", 
"01011011", 
"01111100", 
"10010001", 
"01111000", 
"01010000", 
"10001011", 
"01011011", 
"10001100", 
"10011000", 
"10000010", 
"10010110", 
"01101011", 
"01111001", 
"10000100", 
"01100001", 
"10101001", 
"01110001", 
"00111110", 
"01101110", 
"10011001", 
"01101110", 
"01111110", 
"01111010", 
"01111101", 
"10000101", 
"01011101", 
"10010110", 
"00111111", 
"10010101", 
"10110100", 
"01111010", 
"10010100", 
"01011101", 
"10010010", 
"10011000", 
"01000001", 
"10001101", 
"10101010", 
"10001111", 
"01101111", 
"10001001", 
"01010110", 
"01010011", 
"10100001", 
"10010011", 
"01100000", 
"10010010", 
"01101100", 
"10100001", 
"01010100", 
"01110110", 
"10001011", 
"10011100", 
"01110010", 
"10110010", 
"10010010", 
"01110011", 
"01011111", 
"10001100", 
"01101111", 
"01011101", 
"10000100", 
"01010110", 
"01111001", 
"10001111", 
"10000111", 
"10000001", 
"01011001", 
"10010001", 
"01101000", 
"10000110", 
"10100000", 
"01000111", 
"10010000", 
"10000100", 
"10011101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_0 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_0(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
