use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_81_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_81_LAYER;

architecture Behavioral of ROM_FC_120_81_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_81: ROM_ARRAY_PESOS_FC_120 := (
"01101011", 
"10000000", 
"00111101", 
"10000001", 
"10000000", 
"01000100", 
"10011100", 
"10111000", 
"01110001", 
"01111001", 
"01110110", 
"10001001", 
"01110010", 
"01111000", 
"10001100", 
"10000011", 
"01001111", 
"01101101", 
"10000101", 
"01001110", 
"01111111", 
"00001100", 
"01111001", 
"01110111", 
"01110110", 
"10000100", 
"10000101", 
"01001111", 
"10110100", 
"01010000", 
"10010110", 
"10000010", 
"00101111", 
"01100110", 
"11001001", 
"01000111", 
"10011010", 
"01100100", 
"01001011", 
"01101011", 
"10001010", 
"10101111", 
"10000100", 
"01010100", 
"10101101", 
"00110000", 
"01101010", 
"01110111", 
"01001111", 
"10000000", 
"10000100", 
"10100011", 
"10001110", 
"01110000", 
"00101100", 
"01100100", 
"10001101", 
"10001001", 
"10101000", 
"10011010", 
"01101100", 
"10100101", 
"01100110", 
"01100100", 
"01100011", 
"01111011", 
"01101001", 
"01011001", 
"10010101", 
"10011001", 
"10111110", 
"01100000", 
"01110010", 
"01101100", 
"01100101", 
"01101000", 
"01000000", 
"01110000", 
"01101111", 
"01110001", 
"10001000", 
"10001111", 
"10001000", 
"10011001", 
"01110111", 
"01011000", 
"10001001", 
"01100101", 
"10001000", 
"10001100", 
"01101010", 
"01000101", 
"01100100", 
"01011101", 
"01111111", 
"01100101", 
"10001000", 
"10000111", 
"10001111", 
"01101101", 
"10000101", 
"01111010", 
"10010010", 
"10001001", 
"01110100", 
"01111110", 
"10011100", 
"01101011", 
"01101000", 
"10100001", 
"01110011", 
"10000111", 
"01110111", 
"10110011", 
"01110000", 
"01010110", 
"10000111", 
"01111111", 
"10011010", 
"01001001", 
"10001011", 
"01100111", 
"01011111", 
"10100010", 
"10011000", 
"00110001", 
"01111111", 
"10001100", 
"10001110", 
"10011001", 
"10011010", 
"10000110", 
"10000110", 
"01101111", 
"10010110", 
"01110001", 
"01110010", 
"01101011", 
"10000100", 
"01111001", 
"01101111", 
"10000001", 
"10001000", 
"01110010", 
"10010010", 
"10001011", 
"01101100", 
"10100011", 
"01101110", 
"01111110", 
"01111110", 
"10001000", 
"10001111", 
"01110000", 
"10011010", 
"10001001", 
"10000101", 
"01110001", 
"01110100", 
"01111110", 
"01110110", 
"01100101", 
"10000000", 
"01110110", 
"10010011", 
"10100101", 
"10001110", 
"10111001", 
"10000101", 
"10001000", 
"01111010", 
"10011101", 
"01110110", 
"01100110", 
"10001101", 
"10001000", 
"10011001", 
"01101011", 
"01101011", 
"00010010", 
"01111111", 
"01111110", 
"10001001", 
"10001111", 
"01110111", 
"01110100", 
"01111000", 
"10101111", 
"10000110", 
"01101011", 
"10000001", 
"10001000", 
"10010100", 
"01100110", 
"01110001", 
"10110001", 
"10010110", 
"01101000", 
"01101101", 
"01110110", 
"10000111", 
"10000101", 
"01101001", 
"10000110", 
"01110111", 
"01111101", 
"01110110", 
"01111001", 
"01111101", 
"01101111", 
"01111001", 
"10011111", 
"10001000", 
"10011100", 
"10010101", 
"01010111", 
"01111100", 
"01101101", 
"01110100", 
"10000011", 
"01010111", 
"10110011", 
"10000101", 
"10000100", 
"10100000", 
"01100110", 
"01110110", 
"01010001", 
"01111000", 
"01110001", 
"01111111", 
"10010101", 
"10010001", 
"01110100", 
"10000111", 
"01110101", 
"01110111", 
"01101100", 
"01111100", 
"10001010", 
"01110001", 
"00110010", 
"01110011", 
"01000111", 
"10010101", 
"01010111", 
"10100011", 
"10100010", 
"01110111", 
"10001100", 
"01011101", 
"01110000", 
"01100011", 
"01110010", 
"10000101", 
"01111101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_81: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_81(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
