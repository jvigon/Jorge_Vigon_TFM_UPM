use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_79_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_79_LAYER;

architecture Behavioral of ROM_FC_84_79_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_79: ROM_ARRAY_PESOS_FC_84 := (
"01100011", 
"10001010", 
"10001011", 
"10010110", 
"01100011", 
"10011110", 
"10001111", 
"10000000", 
"10001101", 
"10011101", 
"10001000", 
"01100101", 
"01110110", 
"10001101", 
"01101010", 
"01111111", 
"10001111", 
"01100010", 
"10000111", 
"10001101", 
"01101110", 
"01111101", 
"01011111", 
"01010011", 
"01111011", 
"01011101", 
"10000100", 
"10001010", 
"01110100", 
"10001000", 
"01100101", 
"01010110", 
"01101111", 
"10001101", 
"10011111", 
"01110101", 
"10011110", 
"10001110", 
"01100101", 
"01001001", 
"00011110", 
"10011010", 
"01110011", 
"01110100", 
"01010111", 
"01010101", 
"10000001", 
"01101011", 
"10100110", 
"01101011", 
"01100100", 
"10010010", 
"01110110", 
"01111101", 
"01101001", 
"10000010", 
"10000011", 
"01111100", 
"01011110", 
"10101101", 
"10100001", 
"10100000", 
"10111101", 
"10101100", 
"10100000", 
"10011010", 
"01011110", 
"01110110", 
"10001101", 
"00111100", 
"01100100", 
"01110101", 
"10100110", 
"01101000", 
"10011100", 
"01111000", 
"01100111", 
"10010001", 
"10011101", 
"01000101", 
"01001100", 
"01111100", 
"01010101", 
"01010100", 
"01010010", 
"01110001", 
"10001000", 
"10100010", 
"01101101", 
"01010010", 
"10000000", 
"01111000", 
"10000011", 
"10000001", 
"10110000", 
"01101011", 
"10010000", 
"10000011", 
"01110111", 
"01100000", 
"10011000", 
"01101001", 
"10001001", 
"10010101", 
"01111011", 
"01110110", 
"01101000", 
"10010111", 
"01010000", 
"01101001", 
"01100111", 
"10011001", 
"10000010", 
"11001101", 
"10010000", 
"01101001", 
"10000111", 
"10101100", 
"10001101", 
"01110010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_79: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_79(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
