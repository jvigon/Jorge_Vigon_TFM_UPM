use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_99_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_99_LAYER;

architecture Behavioral of ROM_FC_120_99_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_99: ROM_ARRAY_PESOS_FC_120 := (
"10000010", 
"10010101", 
"01010100", 
"01010011", 
"01110000", 
"10100110", 
"10000110", 
"10000111", 
"10000001", 
"01111110", 
"01111100", 
"10000100", 
"01110001", 
"10010000", 
"01110110", 
"10001101", 
"10001111", 
"10010011", 
"01100111", 
"10001011", 
"01111010", 
"10100011", 
"01111111", 
"01111100", 
"01111001", 
"10000111", 
"01101100", 
"01101011", 
"10010001", 
"01111101", 
"01101110", 
"10001111", 
"10000100", 
"01110111", 
"01111011", 
"10010011", 
"01110000", 
"01111100", 
"10000111", 
"01111100", 
"01110110", 
"01101111", 
"10001011", 
"01110011", 
"01111001", 
"10000000", 
"10010001", 
"01111010", 
"10100000", 
"01101001", 
"10011001", 
"01010000", 
"10001001", 
"01110010", 
"10010101", 
"10011010", 
"10001110", 
"10010100", 
"10000111", 
"01000110", 
"01111101", 
"01101010", 
"01101010", 
"10010000", 
"10001010", 
"01110111", 
"01101101", 
"01101010", 
"01110001", 
"10010001", 
"10110001", 
"01111010", 
"10001000", 
"01100110", 
"01101101", 
"01100000", 
"01000101", 
"01111101", 
"10000000", 
"10001001", 
"10001101", 
"10000101", 
"10001000", 
"10001110", 
"10001001", 
"10110101", 
"01110111", 
"10001000", 
"01111111", 
"01111110", 
"10001110", 
"01110010", 
"01101001", 
"10001110", 
"10001111", 
"01101100", 
"10000100", 
"01100001", 
"10010111", 
"10000110", 
"01110010", 
"01101010", 
"10001000", 
"01011100", 
"01111010", 
"01100001", 
"10011010", 
"01110011", 
"10001000", 
"01011101", 
"01110101", 
"01110000", 
"10010101", 
"10010110", 
"01101111", 
"10100010", 
"01110000", 
"01110011", 
"10010100", 
"01111001", 
"01111010", 
"01111101", 
"10000111", 
"01011100", 
"00111011", 
"10000010", 
"01101100", 
"10001010", 
"10001101", 
"01111000", 
"01111010", 
"01101110", 
"10001000", 
"01110000", 
"01101100", 
"01100111", 
"10001110", 
"01101001", 
"10010010", 
"01111001", 
"10001001", 
"10001100", 
"10001001", 
"10010100", 
"01111111", 
"01101100", 
"01110010", 
"10001010", 
"01111100", 
"01111101", 
"01011001", 
"01111000", 
"10001101", 
"01110100", 
"10000100", 
"10000000", 
"01110010", 
"01101000", 
"01111101", 
"01110011", 
"10010000", 
"01100110", 
"10010100", 
"10100100", 
"10001100", 
"10010000", 
"10000100", 
"10000010", 
"10000010", 
"10010010", 
"10001111", 
"01100101", 
"01101110", 
"01100110", 
"10000000", 
"01101100", 
"01100000", 
"00111111", 
"01110111", 
"10001011", 
"10001011", 
"01100101", 
"01101111", 
"10001111", 
"01110001", 
"10101011", 
"10001110", 
"01110000", 
"01010011", 
"01000101", 
"01101101", 
"10000011", 
"01110001", 
"10010101", 
"00011011", 
"01011000", 
"01101111", 
"10001010", 
"10100101", 
"10000111", 
"10000110", 
"10000100", 
"10000101", 
"10110010", 
"01111001", 
"10000100", 
"10000011", 
"10001010", 
"10010011", 
"01100111", 
"00111100", 
"01011110", 
"01111100", 
"10001000", 
"01111011", 
"10000101", 
"10010000", 
"01011010", 
"01110101", 
"10001111", 
"01000100", 
"01110110", 
"10001110", 
"10001101", 
"01101100", 
"01101100", 
"01110100", 
"01011001", 
"10001101", 
"01010011", 
"01010100", 
"01111001", 
"01111101", 
"01101010", 
"10001100", 
"00111101", 
"00110001", 
"01101110", 
"01110111", 
"10000110", 
"01101100", 
"01011101", 
"01110010", 
"01010111", 
"01111011", 
"01011000", 
"01010111", 
"01110111", 
"01110100", 
"10110001", 
"10001010", 
"01110011", 
"00101100", 
"01011111", 
"10001101", 
"01101111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_99: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_99(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
