use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_58_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_58_LAYER;

architecture Behavioral of ROM_FC_84_58_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_58: ROM_ARRAY_PESOS_FC_84 := (
"01011110", 
"01010001", 
"01110011", 
"10010011", 
"01101011", 
"01110110", 
"10000101", 
"01001101", 
"10111000", 
"10001110", 
"10001010", 
"01111001", 
"10000101", 
"01110110", 
"01111011", 
"01111110", 
"10001100", 
"01100101", 
"01101000", 
"01101011", 
"01110000", 
"01101010", 
"10010101", 
"10101000", 
"01110001", 
"10001100", 
"10011000", 
"01010011", 
"10001100", 
"01111101", 
"10001101", 
"01001011", 
"10000111", 
"10100001", 
"01101110", 
"10011111", 
"10001001", 
"01010110", 
"01100010", 
"01111110", 
"01011100", 
"10010001", 
"01000110", 
"01100111", 
"00101100", 
"01101100", 
"10000001", 
"10010110", 
"01101011", 
"01111000", 
"10011010", 
"00101110", 
"10010001", 
"10011111", 
"01111110", 
"10100100", 
"01100011", 
"10010001", 
"01111000", 
"01101111", 
"01111111", 
"01101101", 
"01010110", 
"01100110", 
"01111010", 
"10011101", 
"01011110", 
"01101110", 
"01111001", 
"01110110", 
"10000101", 
"01010111", 
"10000001", 
"10011000", 
"01110110", 
"10011001", 
"10011011", 
"01111110", 
"01101110", 
"01110001", 
"01100110", 
"01101100", 
"10001000", 
"01100110", 
"01111011", 
"01101110", 
"01011011", 
"10010010", 
"01100011", 
"00111110", 
"10100010", 
"10100101", 
"01111001", 
"00111101", 
"10011010", 
"10011001", 
"10001111", 
"10100100", 
"10100111", 
"01100101", 
"10010110", 
"10000001", 
"01111100", 
"01010101", 
"10001100", 
"10010010", 
"10110010", 
"10001110", 
"00101001", 
"10000110", 
"01000101", 
"01101111", 
"01101100", 
"10010010", 
"01101011", 
"10010111", 
"10010001", 
"10110010", 
"01100101", 
"01101000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_58: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_58(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
