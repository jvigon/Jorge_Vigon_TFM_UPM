use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_33_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_33_LAYER;

architecture Behavioral of ROM_FC_120_33_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_33: ROM_ARRAY_PESOS_FC_120 := (
"10000001", 
"01100100", 
"01101100", 
"01110100", 
"01111001", 
"01100110", 
"01110001", 
"10000100", 
"01110110", 
"10000101", 
"01101111", 
"01011000", 
"01000010", 
"01011001", 
"01101100", 
"10000111", 
"01111110", 
"01000100", 
"01110000", 
"10001101", 
"10000110", 
"10000101", 
"01111110", 
"10001110", 
"01101111", 
"10000001", 
"01111010", 
"01111101", 
"01010101", 
"10001111", 
"10000001", 
"01101100", 
"01101001", 
"01011110", 
"10001001", 
"10100011", 
"10000011", 
"01110100", 
"01011010", 
"10000011", 
"10000110", 
"10000100", 
"01100000", 
"10000110", 
"10000111", 
"01011010", 
"10001001", 
"01111100", 
"01110010", 
"01101100", 
"01110000", 
"01110010", 
"10000101", 
"01111110", 
"01100001", 
"01111100", 
"10000000", 
"01101011", 
"01101010", 
"01111011", 
"01101011", 
"10000100", 
"10001010", 
"10001101", 
"01101111", 
"01100011", 
"10001000", 
"01011101", 
"01111000", 
"01011110", 
"10010010", 
"10001011", 
"01101101", 
"01110111", 
"01101000", 
"10000010", 
"10000101", 
"10001000", 
"10001010", 
"01101111", 
"01110010", 
"10000101", 
"01100111", 
"01110000", 
"10001010", 
"10011001", 
"01011101", 
"01101111", 
"01101000", 
"01111110", 
"10000011", 
"01100100", 
"01101011", 
"01100011", 
"01101010", 
"01110100", 
"01101010", 
"01101011", 
"01101011", 
"10000010", 
"01101111", 
"01010010", 
"01100110", 
"01111000", 
"10000010", 
"10000011", 
"01111011", 
"10001101", 
"01010000", 
"10010000", 
"01101110", 
"10001101", 
"01101100", 
"01100101", 
"01011110", 
"01111111", 
"01110111", 
"01111000", 
"01101100", 
"01101100", 
"01101110", 
"01011100", 
"01101101", 
"10000111", 
"01001110", 
"01110100", 
"01111101", 
"01110010", 
"10001011", 
"10001111", 
"10001111", 
"01011110", 
"10001100", 
"01111110", 
"10100110", 
"01100110", 
"01110000", 
"01101010", 
"10000011", 
"10010101", 
"10010111", 
"01111111", 
"01110011", 
"01110110", 
"10000000", 
"01110001", 
"01111010", 
"01100110", 
"01111010", 
"10001001", 
"01011010", 
"01111011", 
"01110000", 
"01101101", 
"01101101", 
"01100101", 
"01101101", 
"10000001", 
"10001010", 
"01110010", 
"01110110", 
"01001100", 
"01100110", 
"01111101", 
"01111111", 
"01101100", 
"01100010", 
"01101111", 
"01101001", 
"01100101", 
"01101000", 
"01111001", 
"01101001", 
"10011111", 
"10001011", 
"01110000", 
"01111011", 
"01010111", 
"10011000", 
"11100101", 
"10000101", 
"01110011", 
"01111101", 
"01011111", 
"01110110", 
"01100010", 
"01101100", 
"10000110", 
"01101110", 
"10010011", 
"01101010", 
"01110010", 
"01111011", 
"01111100", 
"01010111", 
"01101011", 
"10000010", 
"10000011", 
"01110100", 
"01110110", 
"10000010", 
"01110011", 
"01110111", 
"01010111", 
"01001100", 
"01010110", 
"10001000", 
"10001010", 
"01110000", 
"01101110", 
"01011101", 
"10010011", 
"10000001", 
"01111110", 
"01110110", 
"10000010", 
"10000111", 
"01110100", 
"01101011", 
"10001101", 
"01010101", 
"10001000", 
"10001101", 
"01101001", 
"01111011", 
"10011010", 
"01101110", 
"01100100", 
"10000010", 
"01101110", 
"01111010", 
"10000101", 
"10001011", 
"01011011", 
"01001111", 
"01001110", 
"01111101", 
"10000111", 
"01101010", 
"01111011", 
"01101011", 
"01111010", 
"01110001", 
"10010100", 
"01111101", 
"10000001", 
"10001111", 
"01101111", 
"01111011", 
"01110111", 
"01111101", 
"01101000", 
"01110000", 
"01101111", 
"01111000", 
"01111011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_33: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_33(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
