use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_47_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_47_LAYER;

architecture Behavioral of ROM_FC_120_47_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_47: ROM_ARRAY_PESOS_FC_120 := (
"01110011", 
"01100101", 
"01111000", 
"01100100", 
"01111101", 
"01101001", 
"01010100", 
"01110101", 
"10001101", 
"01110011", 
"01101111", 
"01111001", 
"01001111", 
"01100110", 
"10001010", 
"01110111", 
"01101000", 
"01101010", 
"01011010", 
"01011101", 
"01101011", 
"10011011", 
"01110001", 
"10001011", 
"10000110", 
"01101010", 
"10000001", 
"10001001", 
"01110000", 
"01101100", 
"10001011", 
"01110100", 
"01111000", 
"01011000", 
"01101101", 
"01101101", 
"01111100", 
"01110001", 
"10001010", 
"10001001", 
"01110000", 
"01101110", 
"01011110", 
"10100110", 
"01101111", 
"01110000", 
"10000001", 
"10001001", 
"10000001", 
"01101101", 
"01100000", 
"01001011", 
"01110010", 
"01100011", 
"01111011", 
"01111011", 
"01110000", 
"01100110", 
"01111111", 
"10010110", 
"01000100", 
"01010011", 
"01110001", 
"01111101", 
"01110010", 
"10000011", 
"01110001", 
"01101101", 
"10001000", 
"01111001", 
"01011001", 
"01100111", 
"01110110", 
"01101000", 
"01111101", 
"10001111", 
"10011000", 
"10000100", 
"10001001", 
"01101001", 
"01111100", 
"01111010", 
"01101010", 
"01100001", 
"01101110", 
"10000001", 
"01101011", 
"01110101", 
"10010000", 
"01101110", 
"01101000", 
"01100111", 
"01101101", 
"01101011", 
"10000000", 
"10000111", 
"01111110", 
"01111100", 
"01111101", 
"10001010", 
"10000001", 
"01110001", 
"01110110", 
"10010010", 
"01111000", 
"01101101", 
"10000011", 
"10001100", 
"01110001", 
"10010001", 
"01111011", 
"01110111", 
"01101011", 
"01101010", 
"01011011", 
"10001011", 
"01110000", 
"01011010", 
"01110100", 
"10010011", 
"01110001", 
"01100110", 
"10000001", 
"01110010", 
"01010100", 
"01101010", 
"01110100", 
"10001010", 
"01110010", 
"10001110", 
"01100101", 
"01011001", 
"01100111", 
"01101100", 
"01100001", 
"01110000", 
"01101011", 
"10000100", 
"01011100", 
"10000001", 
"10000001", 
"01100010", 
"01110110", 
"01111100", 
"01101101", 
"10010100", 
"01100111", 
"01100100", 
"10000010", 
"01101011", 
"01011100", 
"01111100", 
"01111101", 
"01101101", 
"01111010", 
"01101110", 
"01111101", 
"01101101", 
"10000011", 
"10001001", 
"01100011", 
"01101001", 
"10010000", 
"01111010", 
"10001110", 
"01111001", 
"10000100", 
"01110001", 
"10000110", 
"01111110", 
"01101101", 
"01010110", 
"01100111", 
"01111001", 
"01101110", 
"10001001", 
"01110000", 
"10001011", 
"01011011", 
"01111111", 
"01110010", 
"01110010", 
"10000000", 
"01111101", 
"10001001", 
"01011011", 
"10000001", 
"01110100", 
"01111001", 
"01111000", 
"01110011", 
"10001000", 
"10000011", 
"01111101", 
"01011100", 
"01011111", 
"01101111", 
"01110010", 
"10001100", 
"01101011", 
"01101011", 
"10000001", 
"10001001", 
"10001110", 
"01100100", 
"01101100", 
"10000111", 
"10001001", 
"01111010", 
"01101011", 
"01110011", 
"10000010", 
"10000100", 
"01011100", 
"01111011", 
"01100101", 
"01101111", 
"01101000", 
"10000111", 
"01110000", 
"01001010", 
"01111110", 
"10000100", 
"01111100", 
"01101101", 
"01111000", 
"01101000", 
"01110111", 
"10001111", 
"01110100", 
"01111111", 
"01110110", 
"10001110", 
"01100001", 
"01111100", 
"01111101", 
"01000010", 
"01101110", 
"01111001", 
"01101110", 
"01110011", 
"01111011", 
"01110100", 
"01100100", 
"01110001", 
"01011110", 
"10011000", 
"10001100", 
"01110101", 
"01100000", 
"01110010", 
"10101001", 
"01110001", 
"01100010", 
"01110110", 
"10001000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_47: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_47(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
