use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_63_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_63_LAYER;

architecture Behavioral of ROM_FC_84_63_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_63: ROM_ARRAY_PESOS_FC_84 := (
"01011101", 
"01100111", 
"01111011", 
"10011000", 
"10110111", 
"01111011", 
"01100100", 
"10011010", 
"10010010", 
"01101111", 
"01101111", 
"01100001", 
"01001111", 
"10001101", 
"10000010", 
"01111111", 
"01011110", 
"01001101", 
"01111011", 
"01100010", 
"10001001", 
"10001011", 
"10010001", 
"01110000", 
"10010100", 
"10100101", 
"01110101", 
"01111100", 
"10010010", 
"10001110", 
"01111000", 
"01110001", 
"01101001", 
"10000000", 
"01011110", 
"01010011", 
"01100111", 
"01101001", 
"01110111", 
"01110010", 
"01110110", 
"11001001", 
"10010011", 
"01100101", 
"01011111", 
"10000111", 
"01111110", 
"01100000", 
"01010100", 
"10000011", 
"01011100", 
"01110110", 
"10001010", 
"01101111", 
"10011010", 
"10100001", 
"10010011", 
"10001001", 
"01110111", 
"01101001", 
"01111101", 
"01110010", 
"10101001", 
"01100101", 
"10000011", 
"01110110", 
"01000110", 
"10011000", 
"01100101", 
"01010010", 
"01110010", 
"01011010", 
"01100001", 
"01101001", 
"10000011", 
"10001101", 
"01110111", 
"10001110", 
"01111101", 
"01101010", 
"10010010", 
"01101110", 
"01011110", 
"01101110", 
"01101101", 
"01101100", 
"01111000", 
"01011101", 
"10001001", 
"01110110", 
"10000001", 
"10100100", 
"01110100", 
"01110110", 
"01110000", 
"10100111", 
"01010010", 
"10011011", 
"01011011", 
"01100001", 
"01110000", 
"10011101", 
"01101100", 
"01100011", 
"01010011", 
"10101101", 
"01110111", 
"10000101", 
"10100010", 
"10100011", 
"10011100", 
"10010111", 
"10001000", 
"01110101", 
"01110011", 
"01110011", 
"01111110", 
"01101101", 
"01111001", 
"10011110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_63 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_63(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
