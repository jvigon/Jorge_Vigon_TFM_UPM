use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_19_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_19_LAYER;

architecture Behavioral of ROM_FC_120_19_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_19: ROM_ARRAY_PESOS_FC_120 := (
"10001010", 
"10101011", 
"01001010", 
"01000100", 
"10000100", 
"01011011", 
"01110001", 
"11000011", 
"10001000", 
"10001001", 
"10100001", 
"10000011", 
"00101000", 
"10000100", 
"10000001", 
"10000101", 
"10011001", 
"10010101", 
"01001101", 
"00111100", 
"01110011", 
"01110000", 
"10001111", 
"10000100", 
"01110100", 
"10011011", 
"01111100", 
"10000111", 
"01001001", 
"01000110", 
"10000001", 
"01111001", 
"10100000", 
"01110110", 
"01110000", 
"01101101", 
"01111001", 
"10100100", 
"01000100", 
"01111001", 
"01111001", 
"01110001", 
"01111010", 
"10011110", 
"00111110", 
"01111100", 
"10000100", 
"01101111", 
"01110000", 
"01011100", 
"01010011", 
"01010110", 
"10000101", 
"01110111", 
"01100110", 
"10011001", 
"10001011", 
"10001011", 
"01111101", 
"01101000", 
"01100001", 
"10000110", 
"01110001", 
"01111100", 
"01110000", 
"01001011", 
"01100010", 
"01010011", 
"01111000", 
"01010100", 
"10011010", 
"10100101", 
"10000101", 
"00101111", 
"01101001", 
"01011110", 
"11000010", 
"01011001", 
"10001000", 
"10010101", 
"11001000", 
"01000110", 
"01110011", 
"10010000", 
"10001000", 
"10010000", 
"10010011", 
"10011011", 
"10000011", 
"01000010", 
"01101101", 
"01100111", 
"10100100", 
"10000110", 
"10000110", 
"01111010", 
"10011110", 
"01011111", 
"01011100", 
"01111101", 
"10001000", 
"01001011", 
"01101000", 
"10011010", 
"01111111", 
"01011000", 
"01101001", 
"01100111", 
"10000100", 
"10000000", 
"10000010", 
"01110110", 
"01110101", 
"10001010", 
"01011100", 
"01101111", 
"01110111", 
"01100101", 
"01010111", 
"10100000", 
"10010010", 
"00110111", 
"01000000", 
"10000101", 
"10100000", 
"10101111", 
"01101010", 
"10010001", 
"01011101", 
"01100100", 
"01111110", 
"01111000", 
"10000111", 
"01011101", 
"10011110", 
"01100110", 
"10001011", 
"10011000", 
"10100000", 
"00011010", 
"01101110", 
"00000110", 
"10001101", 
"10000000", 
"01101001", 
"10001011", 
"10101100", 
"01111100", 
"01110001", 
"01011010", 
"10101000", 
"01100010", 
"01011000", 
"01101111", 
"10101010", 
"01001001", 
"10011011", 
"01011010", 
"01110100", 
"10001101", 
"01010010", 
"11000101", 
"10010010", 
"10011011", 
"01110101", 
"01010001", 
"01010101", 
"01110101", 
"01111100", 
"01010110", 
"10010000", 
"01011000", 
"10100100", 
"10110000", 
"01111001", 
"01111101", 
"01010001", 
"10101110", 
"10000010", 
"10000011", 
"01111000", 
"01110010", 
"10000101", 
"01010100", 
"10000001", 
"01000010", 
"10010110", 
"01010110", 
"10100110", 
"10100010", 
"01111110", 
"01110110", 
"01100101", 
"01011010", 
"00111011", 
"10000101", 
"10001101", 
"01110100", 
"10000100", 
"01111010", 
"10000010", 
"10001101", 
"10001110", 
"00111010", 
"00101010", 
"10000001", 
"01101010", 
"01100111", 
"10000001", 
"01010011", 
"10000111", 
"01110000", 
"01101110", 
"10000100", 
"01110011", 
"01101010", 
"10000001", 
"10010100", 
"10011111", 
"01000110", 
"01010011", 
"01011111", 
"10001010", 
"01111100", 
"01110111", 
"10011000", 
"10001111", 
"10000010", 
"10001011", 
"10011111", 
"01110000", 
"01110111", 
"01110100", 
"01101111", 
"10010110", 
"01011111", 
"10011010", 
"01101100", 
"10001010", 
"10010101", 
"01110010", 
"10001100", 
"01111100", 
"10011010", 
"10000110", 
"01010011", 
"01101011", 
"01100010", 
"01110000", 
"10010100", 
"10001110", 
"10001111", 
"10110000", 
"10000101", 
"10000000", 
"10001000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_19: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_19(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
