LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
use work.CNN_Package_First_Convolution.all;

entity ROM_FIRST_LAYER_POOL is
        Port ( CLK : in STD_LOGIC;
           Reset : in STD_LOGIC;
           addra_pool_1 : IN STD_LOGIC_VECTOR((log2c(Dim_total_Pesos)-1) downto 0);
           douta_pool_1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FIRST_LAYER_POOL;

architecture Behavioral of ROM_FIRST_LAYER_POOL is
SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FIRST is Array (0 to (Dim_total_Pesos-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
CONSTANT ROM_PESOS_FIRST_POOL: ROM_ARRAY_PESOS_FIRST := (
           "10001100", 
        "10010000", 
        "00110000", 
        "10010000", 
        "01011010", 
        "10110010", 
        "00111000", 
        "01101000", 
        "01110011", 
        "10010010", 
        "10110100", 
        "11100011", 
        "11011111", 
        "10100110", 
        "01101001", 
        "01011111", 
        "10001001", 
        "10001111", 
        "01110010", 
        "10000111", 
        "10010111", 
        "00111101", 
        "10001011", 
        "10010011", 
        "10000100", 
        "10100010", 
        "10010100", 
        "10101001", 
        "01110010", 
        "01110100", 
        "01110101", 
        "01011011", 
        "01011110", 
        "10111001", 
        "01110100", 
        "01011000", 
        "10011000", 
        "01100001", 
        "01100000", 
        "10010100", 
        "01111111", 
        "01001001", 
        "01110110", 
        "01100001", 
        "01111101", 
        "10010010", 
        "10011100", 
        "01101111", 
        "01100111", 
        "01000101", 
        "01101111", 
        "10110101", 
        "10001110", 
        "01101010", 
        "10001001", 
        "11001101", 
        "01100100", 
        "00111101", 
        "10100111", 
        "01111011", 
        "10111110", 
        "10001001", 
        "01011101", 
        "01001011", 
        "10110000", 
        "10101000", 
        "01101100", 
        "10001000", 
        "01111111", 
        "01100010", 
        "10110110", 
        "01110100", 
        "01111010", 
        "10000001", 
        "10010110", 
        "10011110", 
        "10010101", 
        "10111011", 
        "10111100", 
        "01011111", 
        "10000010", 
        "01100011", 
        "01010101", 
        "10101110", 
        "10110100", 
        "01101001", 
        "10000010", 
        "01010001", 
        "01010000", 
        "10011110", 
        "01101000", 
        "01101100", 
        "00101111", 
        "01111101", 
        "10100101", 
        "10010111", 
        "10001001", 
        "10010101", 
        "10011101", 
        "10010001", 
        "01110101", 
        "10111010", 
        "10010100", 
        "01111110", 
        "10101010", 
        "10010110", 
        "01100101", 
        "10100110", 
        "01110110", 
        "10001011", 
        "01011010", 
        "10001001", 
        "10001100", 
        "10101000", 
        "10110000", 
        "01010000", 
        "01110000", 
        "01100010", 
        "01011101", 
        "01110010", 
        "10000011", 
        "01100000", 
        "01101110", 
        "01110001", 
        "01100010", 
        "01111011", 
        "10110101", 
        "10100000", 
        "10100001", 
        "01111111", 
        "10100111", 
        "10011010", 
        "01100011", 
        "01111000", 
        "01010101", 
        "10011011", 
        "01100100", 
        "01010111", 
        "01101110", 
        "01011001", 
        "01110000", 
        "01001101", 
        "10000000", 
        "01011101", 
        "10100000", 
        "01010110", 
        "10010010", 
        "10000011", 
        "10010111", 
        "10011010"
);
begin
W_next<= ROM_PESOS_FIRST_POOL(TO_INTEGER(UNSIGNED(addra_pool_1)));
douta_pool_1<= W_reg;
PROCESS (clk,reset)
	BEGIN
		   IF reset='0' THEN
		       
		       W_reg <= (others => '0');
		      
		   elsif CLK'event and CLK='1' then

				W_reg <= W_next;
                      
			END IF;
 end process;

end Behavioral;
