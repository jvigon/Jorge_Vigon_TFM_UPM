use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_94_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_94_LAYER;

architecture Behavioral of ROM_FC_120_94_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_94: ROM_ARRAY_PESOS_FC_120 := (
"01010101", 
"10001000", 
"01111011", 
"01110010", 
"10101111", 
"01101001", 
"01001011", 
"01001001", 
"10000111", 
"01111010", 
"10001100", 
"01110000", 
"10100000", 
"01111101", 
"10010010", 
"01101000", 
"01011010", 
"10001100", 
"01110110", 
"01111001", 
"01111001", 
"01010001", 
"01101010", 
"01101110", 
"01111001", 
"01111111", 
"10001000", 
"10000111", 
"10000010", 
"00111101", 
"01100010", 
"10001001", 
"01011101", 
"01110010", 
"01101101", 
"01111010", 
"01100100", 
"01101010", 
"01111110", 
"10001011", 
"01110101", 
"10000110", 
"10001110", 
"01101101", 
"01101011", 
"01011001", 
"01111111", 
"01011101", 
"10000100", 
"10100110", 
"01100101", 
"10010110", 
"01110111", 
"01110000", 
"01101111", 
"10000011", 
"10000111", 
"10011000", 
"10011010", 
"10101101", 
"01100001", 
"01110110", 
"10010000", 
"01100111", 
"01110101", 
"01100101", 
"01110010", 
"01110101", 
"10011000", 
"00101011", 
"01001010", 
"01110010", 
"01110100", 
"10001100", 
"10010110", 
"10100000", 
"01110111", 
"10100101", 
"01110110", 
"01110110", 
"00110000", 
"01101100", 
"10001100", 
"10010101", 
"01100101", 
"01010111", 
"10011100", 
"10000110", 
"01101010", 
"10000010", 
"01011001", 
"10100000", 
"10100010", 
"01100011", 
"10000101", 
"01100110", 
"01110110", 
"01100100", 
"01101100", 
"01110111", 
"01110100", 
"10001001", 
"01011000", 
"01101011", 
"01101010", 
"10000001", 
"10000100", 
"01101001", 
"10001001", 
"01100001", 
"01100000", 
"10001000", 
"10100001", 
"01111001", 
"01100001", 
"10010011", 
"10000001", 
"01110110", 
"01001000", 
"10100111", 
"01111010", 
"10000100", 
"01110010", 
"01111111", 
"01011011", 
"10000001", 
"10001011", 
"10010101", 
"01110100", 
"01111000", 
"01100010", 
"01010110", 
"01100100", 
"01001110", 
"00111010", 
"01011110", 
"01100100", 
"10001101", 
"01011010", 
"10011010", 
"01110111", 
"11000100", 
"10001101", 
"10010001", 
"01100010", 
"01101010", 
"01000110", 
"01011010", 
"10011101", 
"01001100", 
"01011010", 
"10001100", 
"01111011", 
"10010000", 
"01100000", 
"10011100", 
"01011000", 
"01011101", 
"01111001", 
"01110100", 
"01010011", 
"10001010", 
"01010010", 
"01110001", 
"10001000", 
"10100110", 
"10000110", 
"01110101", 
"01101010", 
"01110011", 
"10100100", 
"10000100", 
"00111011", 
"10001110", 
"01100010", 
"01101100", 
"01110001", 
"11001011", 
"01101110", 
"10100111", 
"10001011", 
"01110101", 
"01110011", 
"01110001", 
"01101101", 
"00011111", 
"01001011", 
"10100000", 
"01101001", 
"10101100", 
"01111110", 
"01110001", 
"10011011", 
"01010101", 
"10011000", 
"01110110", 
"10011100", 
"01010111", 
"10000000", 
"10000001", 
"01111000", 
"01110110", 
"01010110", 
"01111011", 
"10110111", 
"01110111", 
"01110011", 
"10011001", 
"01001111", 
"01111101", 
"10011111", 
"10000001", 
"01110111", 
"00110110", 
"01111001", 
"11011000", 
"01110100", 
"10100010", 
"00101111", 
"01111101", 
"10111111", 
"10100010", 
"10001110", 
"10100000", 
"10010111", 
"10011011", 
"10110110", 
"10100110", 
"10010001", 
"01100111", 
"01111010", 
"10001111", 
"01000101", 
"01111101", 
"01110101", 
"10101100", 
"10001010", 
"10011010", 
"10010110", 
"10001011", 
"10100011", 
"11010110", 
"10001110", 
"01000110", 
"01110000", 
"10011011", 
"01101011", 
"10000010", 
"01101101", 
"01011010", 
"01011110", 
"10010010", 
"11011000", 
"10010110", 
"01110100", 
"10001111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_94: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_94(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
