use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_19_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_19_LAYER;

architecture Behavioral of ROM_FC_84_19_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_19: ROM_ARRAY_PESOS_FC_84 := (
"01011101", 
"01011111", 
"01010101", 
"01111000", 
"01111110", 
"01101100", 
"10001111", 
"01100101", 
"10001001", 
"01001100", 
"10101001", 
"01101010", 
"01110110", 
"10011000", 
"01111101", 
"01110111", 
"10000100", 
"01111111", 
"01011110", 
"01111001", 
"01101111", 
"10100001", 
"10000011", 
"01010100", 
"01111101", 
"10010101", 
"10000001", 
"10001100", 
"01101100", 
"01100101", 
"10010010", 
"10000010", 
"01110010", 
"01111101", 
"10000101", 
"01100100", 
"01100100", 
"01100111", 
"01101111", 
"01101011", 
"01110100", 
"01001101", 
"01011111", 
"10010110", 
"10000001", 
"01100100", 
"01010101", 
"10001111", 
"01011001", 
"01111001", 
"01111001", 
"10000100", 
"01101100", 
"01110100", 
"01111100", 
"10011010", 
"10001110", 
"01110101", 
"10000010", 
"10110110", 
"10000110", 
"01101100", 
"10000011", 
"01010101", 
"01111110", 
"01011000", 
"10101111", 
"10011010", 
"01101001", 
"01111000", 
"10000101", 
"01010100", 
"01110111", 
"01110101", 
"10010010", 
"10011010", 
"10001100", 
"10011101", 
"01111101", 
"01111111", 
"01101100", 
"01010011", 
"01110110", 
"01110100", 
"01101011", 
"10000000", 
"01101101", 
"01101000", 
"01101111", 
"10010001", 
"01110011", 
"01100010", 
"10000100", 
"01111110", 
"01001100", 
"01110010", 
"01111101", 
"01110101", 
"10000100", 
"01110100", 
"10001111", 
"01101100", 
"01110000", 
"01000110", 
"01101000", 
"01101110", 
"10001101", 
"01101001", 
"10000100", 
"10000110", 
"01101111", 
"01101010", 
"10001101", 
"01111001", 
"01110000", 
"10011111", 
"01010101", 
"01111011", 
"10010101", 
"01011001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_19 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_19(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
