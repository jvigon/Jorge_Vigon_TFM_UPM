use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_26_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_26_LAYER;

architecture Behavioral of ROM_FC_84_26_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_26: ROM_ARRAY_PESOS_FC_84 := (
"10001110", 
"10000111", 
"01000100", 
"10010001", 
"01100101", 
"01100110", 
"10001110", 
"01110101", 
"01011110", 
"10000000", 
"01100000", 
"01111111", 
"01110110", 
"10010001", 
"01110101", 
"01111000", 
"01010000", 
"10001011", 
"10010001", 
"01111100", 
"10010110", 
"10000111", 
"10010111", 
"01001111", 
"01111011", 
"01101001", 
"01101000", 
"01111001", 
"00111011", 
"01101000", 
"10000100", 
"00111110", 
"01110001", 
"01101101", 
"01110101", 
"01010010", 
"01011101", 
"10000100", 
"01110001", 
"01101000", 
"01101101", 
"10010000", 
"01010110", 
"01111000", 
"01110010", 
"01111100", 
"01011000", 
"10000011", 
"01101000", 
"01011011", 
"01011111", 
"01010000", 
"10010010", 
"10000011", 
"00101110", 
"01111000", 
"01110110", 
"01100100", 
"10000011", 
"10101111", 
"10001110", 
"01111101", 
"01110011", 
"01000110", 
"01111010", 
"01010010", 
"01101101", 
"10001011", 
"01111101", 
"01111010", 
"01011111", 
"01111011", 
"10001011", 
"01110100", 
"01111000", 
"01111101", 
"11000110", 
"10100001", 
"01101100", 
"01100100", 
"01111110", 
"01110111", 
"01111101", 
"10010001", 
"10101000", 
"10000010", 
"01011011", 
"01101000", 
"10011010", 
"01100100", 
"10101001", 
"10010011", 
"01100110", 
"10011100", 
"10000011", 
"01100111", 
"01100001", 
"10001100", 
"10010010", 
"10001111", 
"10011100", 
"10000000", 
"10001000", 
"01011111", 
"10100010", 
"10000001", 
"10011000", 
"10000011", 
"01001101", 
"10000111", 
"10001111", 
"10000000", 
"01100101", 
"10011100", 
"01110001", 
"01111001", 
"01110011", 
"10111101", 
"10011001", 
"01110011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_26 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_26(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
