use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_22_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_22_LAYER;

architecture Behavioral of ROM_FC_120_22_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_22: ROM_ARRAY_PESOS_FC_120 := (
"10001010", 
"01100011", 
"01010101", 
"01110111", 
"01110001", 
"01111010", 
"01010101", 
"01101100", 
"10000000", 
"01010110", 
"01110110", 
"01111111", 
"01111010", 
"10001000", 
"10001110", 
"10010001", 
"10001001", 
"01001100", 
"01101101", 
"01011011", 
"01011101", 
"10100001", 
"01110101", 
"01101000", 
"10011101", 
"01001100", 
"01111111", 
"01101111", 
"01100011", 
"10100001", 
"01101111", 
"10010011", 
"10011111", 
"01011001", 
"01101100", 
"10100110", 
"10001110", 
"01110101", 
"01110100", 
"01010010", 
"10011110", 
"01100110", 
"01101111", 
"10000101", 
"01111011", 
"01111110", 
"10000000", 
"10000010", 
"01011101", 
"01100001", 
"01111011", 
"01111100", 
"01110011", 
"01100101", 
"01110010", 
"01111000", 
"01111011", 
"01111010", 
"01001110", 
"10000111", 
"01110001", 
"10010110", 
"01110010", 
"01110101", 
"01111101", 
"01100000", 
"01111011", 
"01101110", 
"10000001", 
"01111110", 
"01000011", 
"01111000", 
"10000010", 
"01010100", 
"01101000", 
"01011100", 
"01011110", 
"01111001", 
"01111111", 
"01110101", 
"01111001", 
"01011101", 
"01011010", 
"01001100", 
"10100100", 
"10010001", 
"01111110", 
"01011111", 
"01110101", 
"01111110", 
"01110011", 
"01100001", 
"01101101", 
"10011110", 
"01111011", 
"01110001", 
"01101100", 
"01001111", 
"01101000", 
"10000001", 
"10001101", 
"01100101", 
"01110110", 
"00111101", 
"10011100", 
"01110001", 
"10010111", 
"01101000", 
"01111110", 
"10100001", 
"10001110", 
"10001100", 
"10101010", 
"01101111", 
"01110111", 
"10000000", 
"01110101", 
"01101001", 
"10010101", 
"01010110", 
"10000001", 
"01110111", 
"01001110", 
"10000110", 
"01111000", 
"10000010", 
"10001110", 
"10010010", 
"10001110", 
"10010011", 
"10001001", 
"01101100", 
"01110110", 
"01111000", 
"01011011", 
"10001010", 
"01111010", 
"01101111", 
"01101101", 
"01001110", 
"01101001", 
"10010101", 
"10001000", 
"01111101", 
"10000000", 
"01110010", 
"01011111", 
"01100100", 
"10010101", 
"01110010", 
"10001001", 
"01111010", 
"10011110", 
"01110100", 
"01100011", 
"01101101", 
"01011011", 
"10000001", 
"01111000", 
"01111110", 
"01110001", 
"01101100", 
"01101101", 
"01110001", 
"10000000", 
"01111000", 
"01100000", 
"01000110", 
"01100010", 
"01101101", 
"01101010", 
"10001100", 
"01101101", 
"10100100", 
"01101111", 
"10000000", 
"01110011", 
"01010111", 
"01101010", 
"01101111", 
"01110010", 
"01100001", 
"10100000", 
"01101010", 
"01110010", 
"01111100", 
"01111000", 
"01110111", 
"01110110", 
"01111111", 
"01110101", 
"10000000", 
"10001111", 
"01111001", 
"01011000", 
"01101110", 
"10010011", 
"01011110", 
"01101101", 
"01101011", 
"01111110", 
"01110110", 
"10000101", 
"01111111", 
"01011100", 
"01101001", 
"01110111", 
"10000101", 
"10000100", 
"01011110", 
"01001110", 
"01110110", 
"10001110", 
"01111011", 
"01111100", 
"01100100", 
"10000011", 
"01100111", 
"01011110", 
"01100110", 
"01101111", 
"10000100", 
"10000110", 
"01101101", 
"01100011", 
"01010110", 
"01110011", 
"10000100", 
"10001111", 
"10000000", 
"01111000", 
"01111111", 
"10010101", 
"01101110", 
"01111101", 
"10000100", 
"01101000", 
"01111101", 
"01110111", 
"10000000", 
"10000000", 
"01000111", 
"10000000", 
"01100100", 
"10010010", 
"01011111", 
"01100101", 
"01010100", 
"10001101", 
"01100011", 
"01001111", 
"10000101", 
"01111111", 
"10100100", 
"10000000", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_22: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_22(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
