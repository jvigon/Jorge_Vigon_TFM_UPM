use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_41_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_41_LAYER;

architecture Behavioral of ROM_FC_120_41_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_41: ROM_ARRAY_PESOS_FC_120 := (
"01100101", 
"10111000", 
"10000011", 
"01100100", 
"01110101", 
"01111110", 
"10000110", 
"10001101", 
"10001010", 
"01100100", 
"10010111", 
"10001111", 
"01101001", 
"01101111", 
"10000110", 
"01111000", 
"01100110", 
"00111100", 
"01010011", 
"01111111", 
"01011010", 
"01010100", 
"01010001", 
"01110011", 
"10000110", 
"01010101", 
"10010101", 
"00111100", 
"00110111", 
"01111100", 
"01101111", 
"10000011", 
"01110101", 
"01110000", 
"01100101", 
"11000001", 
"01111011", 
"00111101", 
"01101000", 
"01111110", 
"01110000", 
"01111110", 
"10010001", 
"10010100", 
"01011010", 
"10100000", 
"01101101", 
"10001110", 
"01011001", 
"01101110", 
"01010000", 
"01000010", 
"10000000", 
"01101111", 
"10010000", 
"01100010", 
"10000101", 
"01110101", 
"01110010", 
"01101100", 
"01101000", 
"10000001", 
"01110111", 
"01110001", 
"01100000", 
"01101111", 
"00110011", 
"01111010", 
"01011100", 
"01111111", 
"10001010", 
"01101100", 
"10001110", 
"01001100", 
"01010110", 
"10011001", 
"01100101", 
"01001001", 
"10001011", 
"01110000", 
"10001010", 
"01101110", 
"01100100", 
"01100001", 
"10001101", 
"01100010", 
"01101010", 
"01110010", 
"01111001", 
"01000101", 
"10011010", 
"01010110", 
"01100111", 
"10100001", 
"01111111", 
"01110001", 
"01001110", 
"10000000", 
"01111010", 
"10101000", 
"01110010", 
"01010100", 
"01110110", 
"01000011", 
"01110110", 
"01100100", 
"01110011", 
"10100100", 
"01111010", 
"10011011", 
"10001101", 
"01101100", 
"01010010", 
"10100100", 
"01111000", 
"10010100", 
"10001001", 
"00110011", 
"10000000", 
"00111101", 
"01111011", 
"01111000", 
"01011000", 
"01110000", 
"10011010", 
"10010111", 
"01111011", 
"01110000", 
"01110101", 
"10011000", 
"10000101", 
"00111100", 
"01110101", 
"01011010", 
"01110100", 
"10010100", 
"01111010", 
"01010000", 
"01101110", 
"10001111", 
"01011000", 
"01011000", 
"01101011", 
"10001111", 
"01110000", 
"01010110", 
"10010110", 
"01011010", 
"10000100", 
"01001100", 
"01010111", 
"01110101", 
"10010000", 
"10010001", 
"10000000", 
"01000111", 
"01001100", 
"01000110", 
"01110110", 
"10000010", 
"01100110", 
"01010111", 
"01011111", 
"10010110", 
"01111000", 
"01100001", 
"01001000", 
"01110101", 
"01110010", 
"10010000", 
"10001100", 
"01011001", 
"01101101", 
"01010101", 
"01101100", 
"01111001", 
"01111101", 
"01001111", 
"01100110", 
"10111110", 
"10000000", 
"01111010", 
"01111000", 
"10010100", 
"01111110", 
"10000000", 
"01100000", 
"10100111", 
"01111011", 
"10001011", 
"01101100", 
"01110001", 
"01111111", 
"10000111", 
"10000000", 
"01101101", 
"10000010", 
"01100000", 
"10110011", 
"10000011", 
"10000001", 
"01011111", 
"10011000", 
"10100011", 
"01100000", 
"01001101", 
"10001110", 
"10000101", 
"10000101", 
"01111010", 
"10001100", 
"01101011", 
"01111011", 
"10001101", 
"11000001", 
"10011001", 
"01110010", 
"01111000", 
"10011010", 
"01010010", 
"00110110", 
"01000010", 
"10001101", 
"10001110", 
"01101100", 
"01111101", 
"10010110", 
"01111001", 
"01101100", 
"01011011", 
"01000000", 
"10000010", 
"01111110", 
"01110000", 
"01101110", 
"01100000", 
"00111101", 
"01010100", 
"01111101", 
"01101010", 
"01101100", 
"10000101", 
"01100101", 
"10110000", 
"01111010", 
"01111011", 
"10111010", 
"01000111", 
"01110010", 
"01101001", 
"01110111", 
"01111110", 
"10001000", 
"01100111", 
"10001110", 
"01110000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_41: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_41(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
