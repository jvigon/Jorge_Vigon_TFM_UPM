use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_8_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_8_LAYER;

architecture Behavioral of ROM_FC_120_8_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_8: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"01110011", 
"01000010", 
"01100101", 
"10010000", 
"10100000", 
"10010101", 
"10000100", 
"01110110", 
"01011001", 
"10010111", 
"10110001", 
"10110100", 
"01110001", 
"01110001", 
"01110000", 
"01111000", 
"01010011", 
"10000000", 
"10011101", 
"01111111", 
"10101100", 
"01001010", 
"10010000", 
"10001000", 
"10010101", 
"10101001", 
"01101011", 
"10011011", 
"01101101", 
"01111011", 
"10001000", 
"01110010", 
"01111010", 
"01011011", 
"00110001", 
"01111100", 
"01100001", 
"01111100", 
"01101001", 
"10001110", 
"10100001", 
"01101101", 
"01111011", 
"01110001", 
"10011100", 
"01111110", 
"10001110", 
"01100011", 
"01011110", 
"01101101", 
"10001010", 
"10000101", 
"01111111", 
"10111101", 
"10000110", 
"01111010", 
"01111111", 
"01110001", 
"10000000", 
"11100000", 
"01011001", 
"10010100", 
"10001111", 
"01100101", 
"01000111", 
"01111100", 
"10000011", 
"01111001", 
"10000101", 
"10001110", 
"01110010", 
"10001111", 
"01101011", 
"01111010", 
"01101001", 
"10011010", 
"01011110", 
"01101111", 
"01010100", 
"01110010", 
"01100101", 
"10010100", 
"10011000", 
"10010111", 
"10010010", 
"00110110", 
"01111010", 
"01111110", 
"01111100", 
"10100110", 
"01110000", 
"01001011", 
"01111100", 
"01111100", 
"01101011", 
"01101001", 
"01111110", 
"01101011", 
"01110001", 
"10010001", 
"01011000", 
"01100011", 
"10000010", 
"10000000", 
"01100011", 
"01110110", 
"01100111", 
"10001001", 
"10010001", 
"10010101", 
"01110101", 
"01101110", 
"01111010", 
"01111010", 
"00111100", 
"10000111", 
"01100000", 
"10000011", 
"01111110", 
"01111110", 
"10010110", 
"01110100", 
"10100001", 
"10100001", 
"01100001", 
"10010100", 
"01110001", 
"01100001", 
"01011110", 
"10000000", 
"01011111", 
"01111100", 
"10100011", 
"10010111", 
"01111001", 
"10001011", 
"01100010", 
"10010010", 
"01001100", 
"01100111", 
"01010111", 
"01101111", 
"01110101", 
"01011000", 
"01110101", 
"01111111", 
"10011100", 
"10001111", 
"01100101", 
"01101111", 
"10000111", 
"10000010", 
"10001010", 
"10100111", 
"01111111", 
"01010000", 
"01110101", 
"10000111", 
"01111011", 
"10001101", 
"01001000", 
"01010011", 
"01100001", 
"01111010", 
"01110001", 
"01110011", 
"10010001", 
"01110000", 
"10111000", 
"00110110", 
"01101110", 
"01011110", 
"10001101", 
"10001101", 
"10000000", 
"10000010", 
"01011011", 
"01101001", 
"01111101", 
"10010011", 
"01101100", 
"01101001", 
"10011110", 
"10000111", 
"10101010", 
"01010110", 
"01111010", 
"01101110", 
"01101100", 
"01110101", 
"01110001", 
"10000111", 
"10010111", 
"01111110", 
"01000000", 
"01110110", 
"01101110", 
"10010001", 
"10001101", 
"10001010", 
"01101010", 
"10010111", 
"00100000", 
"10010011", 
"10000100", 
"01101011", 
"01111100", 
"01100110", 
"01010011", 
"01101111", 
"01010110", 
"01111011", 
"11000011", 
"10001110", 
"10011101", 
"01111001", 
"01011100", 
"11000011", 
"01100000", 
"01101100", 
"10100011", 
"01111100", 
"01110010", 
"01011011", 
"01101000", 
"01100010", 
"10010110", 
"01111001", 
"10000010", 
"10111110", 
"01011001", 
"10001001", 
"01110000", 
"10000010", 
"01100000", 
"01101001", 
"10010000", 
"10001010", 
"01101100", 
"01011001", 
"10010111", 
"01111000", 
"10010001", 
"10001111", 
"10000111", 
"01110101", 
"01110000", 
"01111111", 
"01001010", 
"01111011", 
"01111010", 
"01110111", 
"01110110", 
"01110101", 
"01110010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_8 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_8(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
