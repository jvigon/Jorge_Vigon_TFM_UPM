use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_12_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_12_LAYER;

architecture Behavioral of ROM_FC_84_12_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_12: ROM_ARRAY_PESOS_FC_84 := (
"01101011", 
"01100101", 
"10001011", 
"01100100", 
"10000100", 
"01101100", 
"10001000", 
"10100110", 
"01101101", 
"01100000", 
"01110000", 
"01011101", 
"01100010", 
"10010010", 
"10100000", 
"01101010", 
"01000101", 
"01100101", 
"01101011", 
"01100111", 
"10111000", 
"10101001", 
"10001011", 
"10000101", 
"10000010", 
"10100110", 
"01101010", 
"10000100", 
"10001111", 
"10011000", 
"10001111", 
"10001110", 
"10010101", 
"01100010", 
"10000011", 
"01101101", 
"01110001", 
"10001101", 
"10011111", 
"01001010", 
"01100001", 
"10010001", 
"10011000", 
"01101011", 
"01111111", 
"01010100", 
"01100010", 
"10010010", 
"10000001", 
"10010000", 
"10000100", 
"10100100", 
"01110000", 
"01010000", 
"10111001", 
"01111100", 
"01101001", 
"10010001", 
"10001001", 
"01100010", 
"10001011", 
"10110000", 
"01110101", 
"10011011", 
"01111111", 
"01110100", 
"01110101", 
"01111110", 
"10001011", 
"10010000", 
"10000001", 
"10001011", 
"01100001", 
"01111101", 
"10000001", 
"10001111", 
"01111101", 
"01111001", 
"10011101", 
"01111011", 
"10011001", 
"10000110", 
"01100000", 
"10100000", 
"10010001", 
"01001110", 
"01011010", 
"01010101", 
"01011111", 
"01110101", 
"01110011", 
"10011110", 
"10110110", 
"01001011", 
"10011100", 
"10001101", 
"01010101", 
"01110011", 
"01111010", 
"10010001", 
"01111000", 
"10000010", 
"01100010", 
"01110111", 
"01110111", 
"01110101", 
"10101111", 
"10001000", 
"10001011", 
"10100110", 
"01011101", 
"10001100", 
"01111101", 
"10000000", 
"10001110", 
"01110010", 
"10010011", 
"01011101", 
"10001010", 
"01101100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_12 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_12(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
