use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_37_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_37_LAYER;

architecture Behavioral of ROM_FC_84_37_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_37: ROM_ARRAY_PESOS_FC_84 := (
"01001010", 
"01100100", 
"01111001", 
"01110100", 
"10111011", 
"01011111", 
"01111100", 
"01101111", 
"10000011", 
"01110011", 
"01101111", 
"01101011", 
"10000010", 
"10000000", 
"01011111", 
"01100000", 
"01101011", 
"01100110", 
"10000111", 
"01101001", 
"01110100", 
"01111010", 
"01111000", 
"01111111", 
"01110000", 
"10000110", 
"10001110", 
"01100010", 
"01101010", 
"01011101", 
"01101011", 
"01101101", 
"01101111", 
"01100001", 
"01111101", 
"01001110", 
"01110111", 
"01101011", 
"01101100", 
"01101100", 
"01010011", 
"01101011", 
"01111011", 
"01111010", 
"01010011", 
"01110110", 
"01011000", 
"10000101", 
"01011100", 
"10001011", 
"01111010", 
"01110011", 
"10010010", 
"10000010", 
"10010110", 
"01111011", 
"01111001", 
"10001110", 
"01100010", 
"10011001", 
"01111111", 
"01011001", 
"10001001", 
"01010001", 
"01110111", 
"01111010", 
"10011000", 
"10000010", 
"01110111", 
"10011001", 
"01101110", 
"01111110", 
"01100110", 
"01000001", 
"10000101", 
"01111000", 
"10010111", 
"10000111", 
"01110011", 
"10010011", 
"01101100", 
"01110110", 
"01111011", 
"01001101", 
"01101100", 
"01011100", 
"10001000", 
"10000000", 
"01110100", 
"01110011", 
"01100100", 
"10010011", 
"01111101", 
"01101111", 
"01110101", 
"01100010", 
"01100000", 
"10001101", 
"01110011", 
"01101010", 
"10000110", 
"01011010", 
"01110101", 
"01110001", 
"01110101", 
"10001101", 
"01111010", 
"01100110", 
"01110000", 
"10011011", 
"01111000", 
"10001001", 
"10000100", 
"01101001", 
"01110111", 
"01111110", 
"01100011", 
"01101110", 
"10000110", 
"10010001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_37 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_37(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
