use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_42_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_42_LAYER;

architecture Behavioral of ROM_FC_84_42_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_42: ROM_ARRAY_PESOS_FC_84 := (
"01111110", 
"10011110", 
"00010001", 
"10011010", 
"01111000", 
"10000001", 
"10011000", 
"01101100", 
"10001001", 
"10001100", 
"10000001", 
"10010000", 
"10001101", 
"10011000", 
"01111010", 
"10001111", 
"01110100", 
"10101010", 
"01100000", 
"10010101", 
"01101001", 
"10010101", 
"01111001", 
"10100010", 
"01111100", 
"01101010", 
"01111100", 
"01101011", 
"01010100", 
"00111001", 
"01111000", 
"10010100", 
"01110100", 
"10011101", 
"01110101", 
"01010001", 
"10000101", 
"01101000", 
"10101011", 
"11000111", 
"10001000", 
"01001001", 
"01011101", 
"10110101", 
"01111001", 
"10001110", 
"01001100", 
"10010110", 
"01110110", 
"10000110", 
"10101001", 
"01110111", 
"10000100", 
"10001110", 
"10001000", 
"10111001", 
"01011101", 
"10010001", 
"10100100", 
"10001001", 
"10000011", 
"01000101", 
"01111010", 
"01100010", 
"01011001", 
"10000101", 
"10000100", 
"10000111", 
"10000110", 
"10101101", 
"10011010", 
"01111000", 
"01101110", 
"01101001", 
"10010110", 
"01111100", 
"01001110", 
"01110101", 
"01100100", 
"01111100", 
"01011101", 
"01010011", 
"10001110", 
"10010000", 
"01000110", 
"10011110", 
"10000110", 
"01100111", 
"10000000", 
"10100111", 
"01000011", 
"01001110", 
"01101111", 
"01010111", 
"01001001", 
"10001001", 
"01010000", 
"10000111", 
"01110000", 
"10000010", 
"10001001", 
"10010100", 
"01111100", 
"10010100", 
"10001011", 
"10011010", 
"01111010", 
"10001001", 
"10111000", 
"10110010", 
"01111010", 
"01110000", 
"10001000", 
"10000110", 
"01101011", 
"10100000", 
"01110010", 
"00101111", 
"10001001", 
"10011011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_42: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_42(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
