use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_36_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_36_LAYER;

architecture Behavioral of ROM_FC_84_36_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_36: ROM_ARRAY_PESOS_FC_84 := (
"01100110", 
"01111101", 
"10001000", 
"01111001", 
"10101000", 
"10001110", 
"10001111", 
"10000000", 
"01001101", 
"01100101", 
"10001100", 
"01000011", 
"01011100", 
"10100111", 
"01010010", 
"10011111", 
"01010101", 
"01111010", 
"01010011", 
"01101100", 
"10001010", 
"10101100", 
"01110001", 
"01101110", 
"10001011", 
"00110000", 
"01111111", 
"10001100", 
"10000010", 
"10000011", 
"01111011", 
"01101000", 
"10001001", 
"10010001", 
"10001111", 
"01101000", 
"10011111", 
"01110001", 
"10010011", 
"01011100", 
"01011011", 
"11001101", 
"01011011", 
"01101001", 
"10000101", 
"10000011", 
"01010010", 
"10001010", 
"01110100", 
"10010100", 
"10000101", 
"10000101", 
"10001101", 
"01111111", 
"10000001", 
"10001100", 
"01101111", 
"01101011", 
"01100010", 
"01111001", 
"01011100", 
"10001011", 
"01011011", 
"01001110", 
"10011000", 
"01101010", 
"01100110", 
"01110011", 
"10001101", 
"10011110", 
"01110110", 
"01101011", 
"01101110", 
"01111001", 
"10000111", 
"10000100", 
"01100101", 
"01100111", 
"10000011", 
"10000010", 
"01011011", 
"01011011", 
"01111010", 
"01111000", 
"01000101", 
"01111101", 
"10001101", 
"01001001", 
"01110101", 
"01101100", 
"01010111", 
"01101100", 
"10001000", 
"10001100", 
"01101001", 
"01110110", 
"01011100", 
"01110101", 
"01111010", 
"10001010", 
"10011111", 
"10001000", 
"01110010", 
"01011111", 
"01101011", 
"10001001", 
"10010111", 
"01100111", 
"01110001", 
"10110011", 
"10001011", 
"10000110", 
"10010001", 
"10001011", 
"01111101", 
"01101100", 
"10010001", 
"10100101", 
"01110101", 
"10001100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_36 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_36(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
