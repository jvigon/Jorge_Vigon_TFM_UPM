use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_44_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_44_LAYER;

architecture Behavioral of ROM_FC_120_44_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_44: ROM_ARRAY_PESOS_FC_120 := (
"10100101", 
"01101111", 
"01100011", 
"01001111", 
"10011100", 
"01111110", 
"10010111", 
"10011101", 
"01101111", 
"01101111", 
"01110000", 
"01101001", 
"01111010", 
"01110110", 
"01111101", 
"10011100", 
"10001011", 
"10001001", 
"10010011", 
"10010011", 
"10001010", 
"01110110", 
"10001010", 
"01111001", 
"01110010", 
"10010010", 
"01011001", 
"10001001", 
"10000001", 
"01110010", 
"10000110", 
"01101100", 
"10001001", 
"01101001", 
"10101101", 
"01111111", 
"01111100", 
"01111101", 
"10100001", 
"10100011", 
"01111010", 
"01110110", 
"10001011", 
"10000001", 
"10000000", 
"01001010", 
"10000001", 
"10000010", 
"01111000", 
"10001100", 
"01011011", 
"00111100", 
"01111110", 
"01100010", 
"01011000", 
"10011000", 
"01111101", 
"10001000", 
"01101111", 
"01010101", 
"10011111", 
"10000101", 
"01111010", 
"10001010", 
"01101110", 
"01101111", 
"11001001", 
"10110100", 
"01111010", 
"10001000", 
"01101110", 
"01110000", 
"01110100", 
"01111101", 
"01111101", 
"01011100", 
"01100101", 
"10011101", 
"10001110", 
"10001000", 
"10000000", 
"01111011", 
"01110110", 
"10011010", 
"01100010", 
"10001100", 
"01111100", 
"10011100", 
"01111110", 
"10001010", 
"10000000", 
"10010000", 
"01101000", 
"10111111", 
"10010110", 
"10001111", 
"01010100", 
"10010000", 
"10010001", 
"10001110", 
"01101100", 
"10100001", 
"01001011", 
"10000101", 
"10000010", 
"10011000", 
"11010000", 
"10101000", 
"01110110", 
"01010001", 
"10000101", 
"10000100", 
"01110001", 
"10010110", 
"01100011", 
"10010010", 
"01101000", 
"01111000", 
"10011111", 
"01111001", 
"10001110", 
"01011010", 
"10010010", 
"10001100", 
"10010001", 
"01110100", 
"10011100", 
"01011000", 
"10110110", 
"10010110", 
"01111111", 
"10110100", 
"01101111", 
"10001010", 
"01101100", 
"01110010", 
"01110111", 
"10011000", 
"10000101", 
"10000011", 
"01011011", 
"10011111", 
"10000100", 
"01101100", 
"10001001", 
"01101000", 
"01110010", 
"01101011", 
"10001111", 
"01100000", 
"01100111", 
"01111000", 
"01110101", 
"10011100", 
"10011000", 
"10010101", 
"10000011", 
"10101011", 
"10001001", 
"01111001", 
"10010101", 
"10000100", 
"01110100", 
"01010101", 
"10001100", 
"10111101", 
"01010110", 
"10010100", 
"10001000", 
"10010101", 
"10010000", 
"01111000", 
"10011100", 
"00100100", 
"10000001", 
"01110000", 
"01101111", 
"01011100", 
"01100110", 
"01001001", 
"10000100", 
"10010001", 
"10011010", 
"10000000", 
"01110110", 
"10010001", 
"10001110", 
"01110101", 
"01011011", 
"01110101", 
"10011000", 
"01101111", 
"01111000", 
"01100011", 
"00000000", 
"01111011", 
"01111000", 
"11001010", 
"10100111", 
"11000101", 
"01111101", 
"01101011", 
"01110100", 
"10111111", 
"01111101", 
"01011101", 
"01111101", 
"01111001", 
"11110001", 
"01110010", 
"00000000", 
"01001011", 
"10000010", 
"10100011", 
"01111010", 
"10001111", 
"10001001", 
"01001111", 
"01110100", 
"10000001", 
"00110011", 
"01100010", 
"01111100", 
"01100001", 
"10010011", 
"01001111", 
"00111101", 
"01000110", 
"10011110", 
"01101101", 
"01101001", 
"10111101", 
"01111111", 
"10000101", 
"10010110", 
"01011100", 
"00010011", 
"01010101", 
"01101111", 
"01101010", 
"01001110", 
"00000100", 
"10101110", 
"10010101", 
"10000100", 
"01100100", 
"10110100", 
"01110010", 
"10010010", 
"10010001", 
"01111000", 
"01010110", 
"00011111", 
"01101100", 
"10010001", 
"10000110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_44: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_44(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
