use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_20_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_20_LAYER;

architecture Behavioral of ROM_FC_120_20_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_20: ROM_ARRAY_PESOS_FC_120 := (
"01101001", 
"01010100", 
"10100100", 
"10011101", 
"01111011", 
"01111000", 
"10001000", 
"00111001", 
"01110100", 
"10011010", 
"10110101", 
"00111011", 
"10000101", 
"00110111", 
"10001010", 
"01110110", 
"00111000", 
"01111001", 
"10100101", 
"11001001", 
"00110100", 
"01001111", 
"01100001", 
"10011000", 
"01110110", 
"10100110", 
"10011111", 
"01010110", 
"01110001", 
"01010011", 
"01011010", 
"10100111", 
"00101101", 
"01010101", 
"01001111", 
"01100001", 
"01111011", 
"01101000", 
"01001011", 
"10001001", 
"01011011", 
"01110101", 
"01100110", 
"10011101", 
"01001100", 
"01111001", 
"01111111", 
"10001001", 
"01010010", 
"01010010", 
"01010001", 
"10011010", 
"01101110", 
"01101111", 
"00110111", 
"01101000", 
"01110100", 
"01100100", 
"01100001", 
"10100000", 
"01011001", 
"01001000", 
"01011111", 
"01110110", 
"10010011", 
"01100100", 
"10101100", 
"10010000", 
"10111110", 
"10011110", 
"10000011", 
"01000000", 
"10001011", 
"10001110", 
"10100001", 
"01010101", 
"01101000", 
"01011111", 
"01101011", 
"10101011", 
"10010001", 
"10000100", 
"10100010", 
"10010110", 
"10000100", 
"01001100", 
"01010110", 
"10000001", 
"01111101", 
"01111110", 
"10001001", 
"10001001", 
"01111001", 
"10111001", 
"01110110", 
"10101010", 
"01010101", 
"01010111", 
"01101000", 
"00100101", 
"10000111", 
"01101000", 
"01010101", 
"01011000", 
"10000111", 
"01010000", 
"00110101", 
"10100101", 
"10000010", 
"10011100", 
"01101001", 
"01101100", 
"01100011", 
"10000010", 
"01001110", 
"01100001", 
"01110011", 
"01111010", 
"00110100", 
"00111011", 
"01100000", 
"10010111", 
"01010010", 
"10100110", 
"10000111", 
"01111011", 
"01010100", 
"01111100", 
"01011011", 
"01111101", 
"01110111", 
"01000110", 
"01100010", 
"01001001", 
"01010110", 
"10101110", 
"10011101", 
"10001001", 
"01100001", 
"10100110", 
"01110001", 
"01101011", 
"01011101", 
"10001010", 
"01111111", 
"01100010", 
"01110010", 
"01011110", 
"10010001", 
"10010110", 
"00111101", 
"01100001", 
"01110011", 
"10000010", 
"01001101", 
"10001101", 
"10000000", 
"01101110", 
"01111011", 
"01100111", 
"10000100", 
"10000001", 
"01011110", 
"01000101", 
"10001101", 
"01010110", 
"01011011", 
"00111101", 
"01100111", 
"01100000", 
"00110100", 
"01101110", 
"10000100", 
"10111000", 
"10001101", 
"01110000", 
"00111010", 
"10010011", 
"10011000", 
"01111110", 
"10001010", 
"01111111", 
"10101010", 
"01010100", 
"01100110", 
"01110101", 
"01011001", 
"10000001", 
"10000111", 
"01101011", 
"01110010", 
"10000011", 
"10000111", 
"10010011", 
"10001101", 
"01100011", 
"10001010", 
"01101111", 
"10011101", 
"10001000", 
"10000010", 
"01000001", 
"01011010", 
"10101001", 
"01011100", 
"10000101", 
"01101001", 
"10001100", 
"10001100", 
"10000001", 
"01100101", 
"01110110", 
"01100011", 
"01111010", 
"01111101", 
"10100000", 
"01110001", 
"01101110", 
"01100001", 
"01101010", 
"10011110", 
"10000000", 
"01101010", 
"10001001", 
"01111101", 
"10010000", 
"10001100", 
"01001010", 
"01100111", 
"01001110", 
"01111010", 
"01011100", 
"01111101", 
"01001111", 
"01000011", 
"01100111", 
"10111110", 
"10101010", 
"01111011", 
"01100110", 
"01101100", 
"10011010", 
"10010110", 
"01010001", 
"10000011", 
"01101100", 
"10010000", 
"00101111", 
"01101010", 
"10010111", 
"01101110", 
"01110101", 
"10101101", 
"10011001", 
"01110110", 
"10001110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_20: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_20(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
