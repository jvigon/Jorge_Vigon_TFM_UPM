use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_15_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_15_LAYER;

architecture Behavioral of ROM_FC_120_15_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_15: ROM_ARRAY_PESOS_FC_120 := (
"10001010", 
"10001001", 
"10000110", 
"10010110", 
"01110001", 
"10100011", 
"10000100", 
"10000000", 
"10001111", 
"10001101", 
"10100000", 
"01100111", 
"01110100", 
"01111101", 
"01111010", 
"10001010", 
"01111100", 
"10000101", 
"10100101", 
"10101011", 
"01010011", 
"10101110", 
"10100001", 
"01111110", 
"10010100", 
"01110101", 
"10010101", 
"01110100", 
"01111001", 
"10011010", 
"01110011", 
"10100011", 
"01110000", 
"01100011", 
"01111010", 
"10011010", 
"10000111", 
"10100100", 
"01111110", 
"01101101", 
"10001010", 
"01001010", 
"10000011", 
"10001100", 
"01101100", 
"01010100", 
"10001001", 
"01110011", 
"10011010", 
"01101000", 
"10001001", 
"01100100", 
"01101001", 
"01110011", 
"10001101", 
"01110110", 
"10010001", 
"01100111", 
"10000100", 
"10000101", 
"01010111", 
"10001010", 
"10001000", 
"01101110", 
"01100111", 
"01111100", 
"01111000", 
"01100010", 
"10001101", 
"10000001", 
"01111010", 
"01111100", 
"01111101", 
"10011011", 
"01111110", 
"01111000", 
"01101000", 
"01111001", 
"01110011", 
"01111001", 
"01100010", 
"10001101", 
"10000000", 
"10000101", 
"10011100", 
"10001100", 
"01111100", 
"01010011", 
"10001000", 
"10010110", 
"10010110", 
"01111000", 
"10001001", 
"01111100", 
"01111010", 
"01110101", 
"01101001", 
"01000001", 
"10000000", 
"10000010", 
"01110001", 
"10101111", 
"10001110", 
"01111111", 
"10010010", 
"01110001", 
"01110000", 
"01011001", 
"00111100", 
"01110000", 
"01110110", 
"10000110", 
"01100011", 
"01011010", 
"10000011", 
"10011111", 
"10000101", 
"10001100", 
"10010010", 
"10010011", 
"01110111", 
"01110101", 
"01111011", 
"01110011", 
"01101111", 
"10101000", 
"10010101", 
"01110110", 
"01110011", 
"10001000", 
"10000110", 
"01111010", 
"01100101", 
"01111100", 
"01100000", 
"01101101", 
"01111101", 
"01101111", 
"10000011", 
"01110001", 
"10100000", 
"01110110", 
"01111110", 
"10000000", 
"01111110", 
"01010101", 
"10001100", 
"01110010", 
"10001111", 
"10000000", 
"01001011", 
"01100111", 
"10001101", 
"01110110", 
"01111011", 
"01011111", 
"10011100", 
"10010010", 
"01110011", 
"10010000", 
"01101110", 
"01100011", 
"10010011", 
"01111111", 
"01110101", 
"01111110", 
"10000100", 
"01011110", 
"01101101", 
"10001100", 
"01100110", 
"01101001", 
"10000111", 
"01110110", 
"01111110", 
"10000100", 
"01011000", 
"01011000", 
"10000100", 
"10101110", 
"01110011", 
"10110011", 
"10000010", 
"01010101", 
"10010001", 
"01111000", 
"01111001", 
"01101000", 
"01100011", 
"10100011", 
"10001010", 
"10000000", 
"01110101", 
"01111110", 
"01101011", 
"01101110", 
"01111010", 
"10010111", 
"01101101", 
"10000111", 
"10000101", 
"10001000", 
"01101011", 
"01111011", 
"10100101", 
"01100000", 
"10001110", 
"01110010", 
"10000001", 
"01111001", 
"01111000", 
"00111110", 
"01111000", 
"01110001", 
"01100001", 
"01110111", 
"10001010", 
"01101011", 
"01010001", 
"01100001", 
"10001010", 
"01111101", 
"01101100", 
"01111000", 
"10000001", 
"01111011", 
"01011100", 
"01010011", 
"01111111", 
"01111010", 
"10001001", 
"01111110", 
"01110111", 
"01101101", 
"01101111", 
"01110111", 
"10100010", 
"01101000", 
"01110010", 
"01101101", 
"01011011", 
"01100110", 
"01101110", 
"01110011", 
"01101110", 
"10010101", 
"01100001", 
"01001000", 
"01101101", 
"01101000", 
"10111111", 
"10000011", 
"01010011", 
"10010011", 
"10000101", 
"01100110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_15: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_15(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
