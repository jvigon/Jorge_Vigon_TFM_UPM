use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_104_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_104_LAYER;

architecture Behavioral of ROM_FC_120_104_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_104: ROM_ARRAY_PESOS_FC_120 := (
"10000110", 
"01000001", 
"10000011", 
"01000101", 
"01111000", 
"10001110", 
"10010110", 
"01110000", 
"01101001", 
"10011010", 
"01010111", 
"01111001", 
"01110111", 
"01111110", 
"10001010", 
"10101000", 
"10000011", 
"10001001", 
"10000001", 
"01000111", 
"01110110", 
"10010010", 
"01100001", 
"01110011", 
"10000010", 
"01110010", 
"10000000", 
"01011001", 
"01011100", 
"01011110", 
"01101111", 
"10010000", 
"10010010", 
"01010011", 
"10000000", 
"10110010", 
"01110100", 
"01110111", 
"01100000", 
"10011101", 
"10000100", 
"01110001", 
"01101111", 
"10011001", 
"01010101", 
"01010100", 
"10000110", 
"10000110", 
"10001000", 
"01001101", 
"10000110", 
"10111101", 
"01110101", 
"01011010", 
"10000100", 
"10000101", 
"01110100", 
"01101101", 
"01100000", 
"01011111", 
"01111110", 
"10100000", 
"10000100", 
"10100111", 
"10000100", 
"01101111", 
"01010001", 
"01111101", 
"10000010", 
"01011010", 
"01101011", 
"10000111", 
"01110111", 
"01011010", 
"01111111", 
"01110001", 
"01011011", 
"01011000", 
"01110110", 
"01101110", 
"01101010", 
"01100110", 
"10010101", 
"10011001", 
"10001111", 
"01111101", 
"01110011", 
"10011010", 
"10000101", 
"10000101", 
"10001111", 
"01111111", 
"01010000", 
"01110011", 
"10001100", 
"10000010", 
"10000011", 
"01111011", 
"10001000", 
"10000101", 
"10001111", 
"01010111", 
"10000100", 
"01101000", 
"01110011", 
"10101011", 
"01100100", 
"10011111", 
"01110110", 
"10011001", 
"10000100", 
"10000001", 
"01110110", 
"10100011", 
"01111000", 
"10100110", 
"10000011", 
"01101101", 
"01110000", 
"01001111", 
"10001010", 
"01100110", 
"01100111", 
"10001100", 
"10110101", 
"10001000", 
"10000111", 
"10010110", 
"10000001", 
"01111100", 
"10101010", 
"10000111", 
"10000110", 
"01100110", 
"10000111", 
"10010001", 
"10000011", 
"00100111", 
"01101101", 
"01011101", 
"00100001", 
"10000111", 
"10000011", 
"10000001", 
"01101110", 
"01101001", 
"01111010", 
"10000100", 
"01110111", 
"10001100", 
"01111110", 
"01101001", 
"10010000", 
"01011011", 
"01111001", 
"10000010", 
"10000010", 
"10000001", 
"10001010", 
"01110100", 
"01101000", 
"10000100", 
"10110100", 
"10000101", 
"01110010", 
"01000110", 
"10000100", 
"01011100", 
"01110110", 
"10001010", 
"01001010", 
"10001011", 
"10010101", 
"10011010", 
"10000001", 
"10000010", 
"10000011", 
"10101110", 
"10101001", 
"01001000", 
"01110010", 
"01101010", 
"01111011", 
"01100001", 
"01110001", 
"10011101", 
"01100100", 
"01111011", 
"11000101", 
"01101011", 
"10001001", 
"10001101", 
"01101111", 
"10000101", 
"01111110", 
"10000111", 
"10001111", 
"01110100", 
"00101011", 
"01110001", 
"10000001", 
"01111100", 
"01111110", 
"01000000", 
"00000000", 
"10000100", 
"01111000", 
"10000111", 
"01111111", 
"10000010", 
"10000110", 
"01110000", 
"01110000", 
"01111000", 
"01111011", 
"01101000", 
"10010011", 
"01101100", 
"10000001", 
"01010001", 
"00110001", 
"10001001", 
"10001110", 
"01111100", 
"01110010", 
"01000011", 
"10000011", 
"10010000", 
"01111110", 
"10000011", 
"10000100", 
"01110011", 
"10000000", 
"10101111", 
"01011000", 
"10000110", 
"10001010", 
"01110110", 
"10001100", 
"01111010", 
"10010111", 
"01111110", 
"01110100", 
"10000000", 
"10000100", 
"01100011", 
"01011100", 
"10010010", 
"01111011", 
"11000010", 
"01011100", 
"10000010", 
"10100111", 
"01110110", 
"01111110", 
"10010100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_104 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_104(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
