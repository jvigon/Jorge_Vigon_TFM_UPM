use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_73_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_73_LAYER;

architecture Behavioral of ROM_FC_84_73_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_73: ROM_ARRAY_PESOS_FC_84 := (
"10001011", 
"01110000", 
"01110111", 
"10010001", 
"01100001", 
"01110101", 
"01110100", 
"01011111", 
"01100101", 
"01110111", 
"01101111", 
"10011010", 
"01100001", 
"01100011", 
"10000000", 
"10010011", 
"01011111", 
"10001010", 
"10001110", 
"01111110", 
"01101110", 
"10000011", 
"01100001", 
"01110001", 
"10010100", 
"10010010", 
"10001101", 
"01011111", 
"01110000", 
"10010110", 
"10010010", 
"10010111", 
"01100111", 
"01110100", 
"10001101", 
"01100111", 
"01010100", 
"01111101", 
"01110100", 
"10110111", 
"01110111", 
"10011101", 
"10001010", 
"01000010", 
"01100101", 
"10000110", 
"01011001", 
"01101100", 
"01011111", 
"01101101", 
"10000011", 
"01111111", 
"10000011", 
"01000101", 
"01011101", 
"01100101", 
"01111011", 
"10001001", 
"01110111", 
"10010001", 
"10000100", 
"01010110", 
"10001110", 
"01101100", 
"10000100", 
"01100101", 
"01110100", 
"10000101", 
"10010111", 
"01110010", 
"01111011", 
"10001100", 
"01010100", 
"01100101", 
"01101110", 
"10000110", 
"10010110", 
"01100100", 
"01011100", 
"10001100", 
"01011100", 
"01010010", 
"01100100", 
"10000001", 
"00110101", 
"01110010", 
"10000001", 
"01011101", 
"10010110", 
"01101010", 
"01010001", 
"10001110", 
"01110111", 
"01000110", 
"01110111", 
"10001101", 
"01011001", 
"10011001", 
"01101111", 
"01110101", 
"01101000", 
"10100111", 
"01101101", 
"01100101", 
"01010110", 
"01100110", 
"10010001", 
"01100100", 
"01101010", 
"01101111", 
"01111010", 
"01110111", 
"10000011", 
"10010100", 
"01100101", 
"01110110", 
"01100100", 
"01100111", 
"10001101", 
"01101110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_73: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_73(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
