use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_16_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_16_LAYER;

architecture Behavioral of ROM_FC_84_16_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_16: ROM_ARRAY_PESOS_FC_84 := (
"10100000", 
"10101001", 
"10010001", 
"01111101", 
"10011110", 
"01101001", 
"01110100", 
"01011000", 
"10000001", 
"10010000", 
"10010010", 
"01111010", 
"10000010", 
"10011100", 
"10110101", 
"10001011", 
"01111101", 
"01111010", 
"10101100", 
"10000111", 
"01110110", 
"01010110", 
"01101110", 
"01111011", 
"01100110", 
"10110011", 
"01101100", 
"01011101", 
"10001110", 
"01110000", 
"10001110", 
"10010011", 
"01001110", 
"10010101", 
"01011111", 
"01101001", 
"10100000", 
"01100001", 
"01011010", 
"01101111", 
"01011111", 
"01010110", 
"01110101", 
"00110111", 
"10000101", 
"10100000", 
"10000100", 
"01101000", 
"10100010", 
"10000100", 
"01011100", 
"10100101", 
"10001011", 
"10000111", 
"01010111", 
"10100011", 
"01110111", 
"01100001", 
"01010111", 
"10000001", 
"10100000", 
"01101110", 
"01111100", 
"01111100", 
"10010011", 
"01001111", 
"01011111", 
"01110000", 
"10000000", 
"01010101", 
"10010101", 
"10011101", 
"10010011", 
"01011111", 
"10011000", 
"10001010", 
"01111010", 
"01101101", 
"10011000", 
"10001000", 
"10001001", 
"01111010", 
"01101000", 
"01100000", 
"01101111", 
"01101101", 
"10011000", 
"10110000", 
"10001100", 
"10110110", 
"01001111", 
"10100010", 
"10001001", 
"10000100", 
"01101101", 
"10001110", 
"10011011", 
"01101110", 
"01001111", 
"01110010", 
"10001100", 
"01111010", 
"01001100", 
"01010010", 
"10011101", 
"01010111", 
"01000100", 
"10001011", 
"10011000", 
"01001001", 
"01101101", 
"10001010", 
"01110100", 
"10011000", 
"01101100", 
"10000011", 
"01101000", 
"01110011", 
"10011010", 
"01011100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_16 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_16(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
