use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_23_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_23_LAYER;

architecture Behavioral of ROM_FC_84_23_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_23: ROM_ARRAY_PESOS_FC_84 := (
"01011000", 
"01100100", 
"01100111", 
"01110000", 
"10101001", 
"01100010", 
"10001001", 
"01010111", 
"01111110", 
"10010101", 
"10011101", 
"10001110", 
"01001001", 
"01011011", 
"10001001", 
"01001011", 
"01100111", 
"10000101", 
"01011001", 
"01110000", 
"10000101", 
"01101011", 
"01101110", 
"00110100", 
"10000100", 
"10010110", 
"10001110", 
"01011001", 
"01111110", 
"01101011", 
"01111101", 
"10011011", 
"01111010", 
"10000011", 
"00111100", 
"10010000", 
"10011000", 
"01100101", 
"01101101", 
"01100111", 
"01101110", 
"10100000", 
"10000000", 
"01001100", 
"01001010", 
"01111110", 
"11010011", 
"01111101", 
"10001001", 
"01110011", 
"01100111", 
"10110110", 
"10001010", 
"10100110", 
"01110011", 
"10100100", 
"01110000", 
"10010110", 
"01111100", 
"01100110", 
"01111010", 
"01111111", 
"10101001", 
"01110001", 
"10110011", 
"01000100", 
"10011110", 
"01100111", 
"10010001", 
"10001111", 
"10000010", 
"01000101", 
"00111011", 
"01110010", 
"01101111", 
"10001110", 
"01011111", 
"10011001", 
"01101110", 
"10111000", 
"01010101", 
"10011100", 
"00110111", 
"01101101", 
"01110110", 
"01011101", 
"10011010", 
"00111011", 
"10001011", 
"10100111", 
"01111010", 
"01110001", 
"10010010", 
"10011110", 
"01100011", 
"10001000", 
"10010000", 
"10000011", 
"01011110", 
"01010001", 
"01101000", 
"10000010", 
"01101011", 
"01101011", 
"01010111", 
"10010110", 
"01111100", 
"10010001", 
"10010011", 
"10100100", 
"10000001", 
"01111001", 
"01100101", 
"10001010", 
"01110100", 
"10111101", 
"10001000", 
"01001111", 
"01111110", 
"01001010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_23 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_23(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
