use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_72_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_72_LAYER;

architecture Behavioral of ROM_FC_120_72_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_72: ROM_ARRAY_PESOS_FC_120 := (
"01111100", 
"01100100", 
"01111011", 
"10000100", 
"01111010", 
"10110100", 
"10011101", 
"01101010", 
"10000100", 
"01010110", 
"10011110", 
"00001110", 
"10011001", 
"00111110", 
"01111111", 
"10001110", 
"10010111", 
"01011100", 
"10010010", 
"10001010", 
"10100001", 
"10111101", 
"01100011", 
"01111110", 
"01111011", 
"01100010", 
"01101000", 
"01001111", 
"01111111", 
"01110110", 
"10001000", 
"01111111", 
"10110100", 
"01101001", 
"10100001", 
"10001111", 
"10100101", 
"01100100", 
"10001010", 
"10010100", 
"01111111", 
"10001010", 
"10000000", 
"01101110", 
"01110010", 
"01101101", 
"01101001", 
"01110000", 
"10000110", 
"10100011", 
"10100000", 
"01110110", 
"01110100", 
"01100110", 
"01111001", 
"10111110", 
"01100011", 
"10001011", 
"01001101", 
"10000111", 
"01011100", 
"01101000", 
"01101100", 
"01100011", 
"01111000", 
"10101110", 
"01011101", 
"10000100", 
"01111100", 
"01011010", 
"10011011", 
"10000110", 
"10001111", 
"01010011", 
"01110001", 
"10000001", 
"10010000", 
"01000100", 
"10001100", 
"01111000", 
"01100111", 
"01001111", 
"10010000", 
"10011100", 
"10000000", 
"01111010", 
"10111110", 
"10011001", 
"01101010", 
"01010100", 
"10001001", 
"01011110", 
"10001011", 
"10001010", 
"10011010", 
"01101111", 
"10100000", 
"01110101", 
"10000100", 
"01111011", 
"10010100", 
"01101010", 
"01111110", 
"10000100", 
"10000111", 
"10010011", 
"01110101", 
"01100110", 
"10000110", 
"10100001", 
"10000011", 
"01101011", 
"10001010", 
"10011100", 
"10010101", 
"01100000", 
"10000000", 
"01001111", 
"01000001", 
"10101010", 
"10000110", 
"10100100", 
"00100010", 
"10000011", 
"10110110", 
"01110111", 
"01011001", 
"10000101", 
"01111100", 
"10100011", 
"01100000", 
"01101101", 
"10101001", 
"10001011", 
"11001111", 
"01110100", 
"01101110", 
"01000100", 
"01110110", 
"10101101", 
"11000110", 
"00000111", 
"10001010", 
"10000111", 
"01010010", 
"10010110", 
"10001001", 
"10001001", 
"01110111", 
"01011011", 
"10001101", 
"10001001", 
"01110001", 
"01110000", 
"10010100", 
"01011111", 
"10010001", 
"00011111", 
"01100110", 
"10010010", 
"01100011", 
"01100101", 
"10000011", 
"10001100", 
"10000100", 
"10010000", 
"01111000", 
"10010100", 
"10001100", 
"10001011", 
"10101000", 
"10001100", 
"10000001", 
"10001110", 
"01100011", 
"01101010", 
"01011111", 
"10111011", 
"10010000", 
"01111010", 
"10001110", 
"01110111", 
"00111101", 
"10100100", 
"10000110", 
"01101111", 
"01011111", 
"10000010", 
"01010000", 
"10010101", 
"01111110", 
"01111000", 
"10010110", 
"10001011", 
"01111111", 
"10011000", 
"11000100", 
"00100010", 
"01001111", 
"00100010", 
"10001010", 
"01111001", 
"01100001", 
"01100001", 
"01010000", 
"00101010", 
"10000100", 
"01111101", 
"00100111", 
"01100010", 
"10000110", 
"10100000", 
"10001011", 
"10010101", 
"01101111", 
"01001011", 
"01111110", 
"10011100", 
"10011101", 
"00001000", 
"01101001", 
"01010111", 
"01110010", 
"10011010", 
"01100010", 
"01100011", 
"10010001", 
"01111101", 
"10010001", 
"10000010", 
"01001101", 
"01101011", 
"10000010", 
"01111100", 
"10010011", 
"01101110", 
"01100101", 
"01110010", 
"01111101", 
"10000111", 
"10011111", 
"10100101", 
"01111100", 
"01010110", 
"10001110", 
"10010110", 
"10110111", 
"01101101", 
"01111110", 
"01101100", 
"01011011", 
"10001011", 
"10101100", 
"10110100", 
"01100100", 
"10011001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_72: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_72(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
