use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_42_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_42_LAYER;

architecture Behavioral of ROM_FC_120_42_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_42: ROM_ARRAY_PESOS_FC_120 := (
"10001101", 
"10000111", 
"01111011", 
"01000110", 
"10001010", 
"01100100", 
"01110001", 
"01100111", 
"01101011", 
"01011100", 
"01100110", 
"10010011", 
"01111000", 
"01101011", 
"01101010", 
"10001111", 
"10000101", 
"01100111", 
"10010110", 
"01000100", 
"01100101", 
"01001111", 
"01110111", 
"01001000", 
"01110111", 
"01011001", 
"10001010", 
"10001011", 
"10001000", 
"01111111", 
"01111111", 
"10001111", 
"01001111", 
"10001010", 
"01011000", 
"01011111", 
"10000100", 
"01101101", 
"01011001", 
"01111011", 
"10001000", 
"10000011", 
"10101000", 
"01100100", 
"01110011", 
"01101011", 
"01111011", 
"01111010", 
"01110011", 
"01100111", 
"01101011", 
"10010101", 
"10001110", 
"01111000", 
"01101110", 
"10000000", 
"01101001", 
"10001011", 
"10110111", 
"01101010", 
"01100011", 
"01110000", 
"01101110", 
"10001100", 
"01110101", 
"01100110", 
"01110010", 
"10001100", 
"01111001", 
"10000110", 
"00111101", 
"01100101", 
"01110111", 
"01010111", 
"01110011", 
"01100101", 
"01110101", 
"10010110", 
"01101010", 
"10001010", 
"10010010", 
"10001111", 
"01111000", 
"10001001", 
"01101000", 
"01101001", 
"00010001", 
"01011110", 
"01111011", 
"01011010", 
"01111011", 
"01101000", 
"00101010", 
"01110111", 
"01111100", 
"01110101", 
"01100010", 
"10010111", 
"01110110", 
"01001101", 
"01101111", 
"01110000", 
"01111101", 
"01011110", 
"01111010", 
"01011110", 
"10001000", 
"01111100", 
"01001110", 
"10001001", 
"01111110", 
"01110000", 
"01101111", 
"01111000", 
"01011110", 
"10111010", 
"10000100", 
"10010100", 
"10010100", 
"01001000", 
"01101010", 
"00110000", 
"10001110", 
"10000111", 
"00111001", 
"01100011", 
"10010000", 
"01110101", 
"01101011", 
"01010010", 
"10011010", 
"10001111", 
"01110001", 
"01110110", 
"00110010", 
"01011010", 
"01110000", 
"00111100", 
"10011111", 
"01000011", 
"01111101", 
"10100110", 
"01101111", 
"10000001", 
"01100100", 
"01100011", 
"10000100", 
"10001010", 
"10000110", 
"10001110", 
"01111001", 
"10000010", 
"10011100", 
"01101111", 
"01010010", 
"01000111", 
"01100111", 
"10100110", 
"10001001", 
"01111100", 
"01100110", 
"01100010", 
"10001101", 
"10001000", 
"10000010", 
"01110101", 
"11000001", 
"01111011", 
"10000101", 
"01010111", 
"01110000", 
"10100011", 
"01110001", 
"10000100", 
"01110001", 
"01111100", 
"01111111", 
"01101111", 
"01010101", 
"01100010", 
"01111011", 
"01111101", 
"10101111", 
"01010000", 
"10000011", 
"01100000", 
"10001110", 
"01110011", 
"10000110", 
"00111110", 
"01111001", 
"01111101", 
"01110101", 
"01010001", 
"10001001", 
"10000000", 
"10001110", 
"10010001", 
"01010110", 
"01011100", 
"01110001", 
"01111100", 
"10010101", 
"00111100", 
"01100100", 
"01110001", 
"10000010", 
"01111011", 
"01111111", 
"01001101", 
"01100001", 
"10011100", 
"10000010", 
"00111100", 
"01111100", 
"01100110", 
"01110111", 
"01110100", 
"01100101", 
"00000000", 
"01100010", 
"10111111", 
"01111010", 
"01110010", 
"01101010", 
"01100110", 
"10011000", 
"10111100", 
"01111110", 
"01100000", 
"10100010", 
"01010001", 
"01101100", 
"10000000", 
"01100000", 
"00111010", 
"10011011", 
"01100101", 
"10000000", 
"10010011", 
"10011110", 
"10000011", 
"01111001", 
"01100100", 
"01111100", 
"01101101", 
"01110100", 
"10001001", 
"01111011", 
"10101011", 
"10000001", 
"01001001", 
"01110101", 
"01101111", 
"01101011", 
"10001010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_42: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_42(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
