use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_34_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_34_LAYER;

architecture Behavioral of ROM_FC_120_34_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_34: ROM_ARRAY_PESOS_FC_120 := (
"01011000", 
"01110001", 
"10001001", 
"01010000", 
"10011000", 
"00110100", 
"00011000", 
"00111101", 
"10000101", 
"10001110", 
"01111011", 
"11011101", 
"10110111", 
"01110011", 
"01111001", 
"01101110", 
"01011111", 
"10000111", 
"01110100", 
"01110000", 
"01010001", 
"10010101", 
"00100100", 
"01010000", 
"01101110", 
"01000011", 
"01000100", 
"11110001", 
"10100011", 
"10100100", 
"10001100", 
"01111110", 
"10110111", 
"10001100", 
"01000010", 
"01011100", 
"01110111", 
"10101011", 
"01111110", 
"10010010", 
"01111101", 
"01001100", 
"01101010", 
"10010111", 
"01111010", 
"10010000", 
"10001111", 
"10000000", 
"11000100", 
"10010111", 
"10000010", 
"10011111", 
"01110101", 
"01111110", 
"10111000", 
"01011000", 
"01101101", 
"01010110", 
"10100010", 
"00011110", 
"01101100", 
"10001001", 
"10001100", 
"10000101", 
"01110001", 
"01110010", 
"01011000", 
"01011110", 
"01111011", 
"10000001", 
"00110101", 
"01110011", 
"01110111", 
"10000111", 
"01101010", 
"11001010", 
"10000111", 
"10111000", 
"10001111", 
"01111011", 
"01001001", 
"01101111", 
"01011101", 
"01100000", 
"10000011", 
"01111010", 
"01011110", 
"01110111", 
"01111110", 
"10001001", 
"01001011", 
"10000110", 
"10010001", 
"01010110", 
"01111000", 
"10000110", 
"01101010", 
"01010110", 
"10000001", 
"01111110", 
"01110001", 
"01101100", 
"01010010", 
"10101000", 
"01011101", 
"10010111", 
"10000001", 
"01000011", 
"01111101", 
"00011000", 
"01110011", 
"10000011", 
"01100001", 
"00110011", 
"10011111", 
"10110011", 
"01101110", 
"01011101", 
"01100010", 
"10101010", 
"01011100", 
"01100010", 
"01111110", 
"01001101", 
"00011011", 
"10001000", 
"10001001", 
"10001011", 
"10110110", 
"00100011", 
"01011011", 
"01011011", 
"01000001", 
"10010100", 
"00010000", 
"01000100", 
"01111100", 
"01100001", 
"00110001", 
"01110110", 
"01100000", 
"10111111", 
"10001000", 
"01111111", 
"01011111", 
"01110101", 
"01010011", 
"01001011", 
"10010100", 
"01110001", 
"10000110", 
"10100000", 
"01101010", 
"01111111", 
"00100010", 
"10001100", 
"01101001", 
"10011100", 
"10010010", 
"10001010", 
"01110000", 
"10010100", 
"01011100", 
"01101111", 
"01111001", 
"01110101", 
"10010000", 
"10000010", 
"01100110", 
"10001111", 
"01110101", 
"10010011", 
"01011111", 
"01001111", 
"01100101", 
"10001011", 
"01110101", 
"10010001", 
"10010001", 
"10001011", 
"10000110", 
"01100110", 
"01101000", 
"01001111", 
"01111100", 
"01101101", 
"01100010", 
"10000011", 
"01101010", 
"10011101", 
"10000111", 
"01110001", 
"01111001", 
"00100001", 
"10100111", 
"01110110", 
"01011100", 
"10001101", 
"01011111", 
"10001101", 
"01110011", 
"01111110", 
"01110010", 
"01110101", 
"10101000", 
"01110101", 
"01111011", 
"10000111", 
"01010101", 
"01010100", 
"10000010", 
"01100101", 
"01110110", 
"01001110", 
"11001101", 
"10001001", 
"01111111", 
"01111101", 
"01011000", 
"10011001", 
"10011100", 
"10100111", 
"01111111", 
"10010001", 
"10100101", 
"10010101", 
"01101110", 
"01000110", 
"01101111", 
"01010111", 
"10011100", 
"10000100", 
"01110011", 
"01110010", 
"00101111", 
"10101000", 
"10010111", 
"10001111", 
"01110000", 
"10000100", 
"10011100", 
"10001010", 
"01011000", 
"00100010", 
"01110010", 
"10010011", 
"01101001", 
"10000010", 
"10000110", 
"01111101", 
"01011011", 
"01111000", 
"10101001", 
"01101111", 
"10000000", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_34: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_34(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
