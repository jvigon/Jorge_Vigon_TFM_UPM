use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_3_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_3_LAYER;

architecture Behavioral of ROM_FC_84_3_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_3: ROM_ARRAY_PESOS_FC_84 := (
"01101010", 
"10000100", 
"10000100", 
"01110000", 
"10000000", 
"01101111", 
"10010101", 
"01101001", 
"10000111", 
"01101000", 
"01111101", 
"01110101", 
"01101110", 
"10000111", 
"01111110", 
"01001101", 
"01011110", 
"10100000", 
"10010010", 
"01011101", 
"10011101", 
"10000011", 
"10001100", 
"10000110", 
"10000001", 
"10010011", 
"01111100", 
"01011001", 
"01111011", 
"01100101", 
"10001100", 
"01011000", 
"01100001", 
"10010100", 
"10010000", 
"01100100", 
"10101010", 
"01111001", 
"10001010", 
"01011111", 
"10001000", 
"01101110", 
"01110000", 
"01011000", 
"01011110", 
"01111000", 
"01100011", 
"01100110", 
"01111001", 
"01111111", 
"10000110", 
"01111000", 
"10001011", 
"01110100", 
"01111010", 
"01111101", 
"10000100", 
"01101100", 
"01110010", 
"01101000", 
"01111100", 
"10000111", 
"01111111", 
"01011100", 
"10001101", 
"01110011", 
"01101011", 
"01111111", 
"10011001", 
"10010011", 
"01101101", 
"01010101", 
"01100010", 
"01101101", 
"10001001", 
"10000110", 
"10011100", 
"01101110", 
"10000011", 
"01100001", 
"01100001", 
"01111010", 
"01011101", 
"01101101", 
"01100101", 
"10000101", 
"01011101", 
"01111101", 
"01110001", 
"10001000", 
"01110100", 
"10001110", 
"10001100", 
"10000001", 
"01010100", 
"10011000", 
"01001111", 
"10010001", 
"10000001", 
"01011110", 
"10001101", 
"01111100", 
"01110001", 
"01101110", 
"01110101", 
"10010101", 
"10010011", 
"10001000", 
"01010111", 
"10011011", 
"01101011", 
"10010101", 
"01101111", 
"10000000", 
"10011010", 
"01100010", 
"10000010", 
"01110011", 
"01101001", 
"01011010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_3 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_3(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
