use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_7_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_7_LAYER;

architecture Behavioral of ROM_FC_120_7_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_7: ROM_ARRAY_PESOS_FC_120 := (
"01001100", 
"10010010", 
"10011010", 
"01011000", 
"01011010", 
"01101101", 
"01100101", 
"00101111", 
"10010001", 
"10000101", 
"01011011", 
"10100001", 
"01110101", 
"01100001", 
"10000101", 
"01100101", 
"01100010", 
"01111110", 
"10000010", 
"10111001", 
"10000110", 
"10011000", 
"01110000", 
"01100001", 
"01111000", 
"01110111", 
"11000101", 
"10100011", 
"10001010", 
"10010001", 
"01101000", 
"10000011", 
"01110111", 
"01111000", 
"10001011", 
"10100110", 
"01101101", 
"01111001", 
"01110001", 
"10010000", 
"10011100", 
"10011001", 
"10011001", 
"01100010", 
"01011101", 
"01100011", 
"10000001", 
"01110000", 
"01011101", 
"01001100", 
"01101000", 
"01100010", 
"10001000", 
"01011000", 
"10000111", 
"10000100", 
"01111010", 
"10110110", 
"01111000", 
"10010101", 
"01111001", 
"00101001", 
"10000110", 
"10000110", 
"10001111", 
"01101101", 
"01101000", 
"01101111", 
"01010000", 
"00110110", 
"01011000", 
"00110001", 
"10001100", 
"10101100", 
"01111111", 
"10100000", 
"01000010", 
"11000010", 
"10000110", 
"10010000", 
"10011111", 
"01110110", 
"01110110", 
"01111100", 
"01101110", 
"01101001", 
"00101101", 
"01100110", 
"10000101", 
"10010101", 
"10110000", 
"10000111", 
"01100011", 
"10010010", 
"10100000", 
"01101011", 
"01011111", 
"01101000", 
"01100110", 
"01101101", 
"10001100", 
"10011110", 
"00110101", 
"01100001", 
"10001111", 
"01111010", 
"10001001", 
"01000110", 
"01010101", 
"10110000", 
"10000010", 
"01111010", 
"01001011", 
"01000001", 
"01110101", 
"01001100", 
"10010011", 
"01111110", 
"01111011", 
"01110011", 
"10000000", 
"10000010", 
"01011000", 
"10110000", 
"10100011", 
"10101111", 
"10010000", 
"01111000", 
"10011001", 
"01100001", 
"10110000", 
"01011101", 
"01001001", 
"01001101", 
"00110010", 
"10010011", 
"01111101", 
"10110111", 
"01001101", 
"01111001", 
"10001110", 
"10000100", 
"10000011", 
"10010101", 
"01100100", 
"01100001", 
"10001001", 
"01101110", 
"01101111", 
"01111110", 
"01010010", 
"10100011", 
"01110111", 
"10010010", 
"01011111", 
"10011010", 
"01011111", 
"10011101", 
"10000000", 
"01101101", 
"10011001", 
"10000100", 
"01110101", 
"01111011", 
"01110101", 
"10100000", 
"01111000", 
"01100100", 
"10010111", 
"01110011", 
"01110010", 
"10010100", 
"01101101", 
"10110110", 
"10001001", 
"01110111", 
"10000111", 
"10100011", 
"10011111", 
"10100000", 
"10001101", 
"10001010", 
"10011111", 
"01101001", 
"10001111", 
"01001101", 
"01001011", 
"10001001", 
"10100111", 
"10100110", 
"01100101", 
"01111101", 
"10101001", 
"01100011", 
"10010010", 
"01010011", 
"01100100", 
"01100111", 
"10101000", 
"11000110", 
"10000011", 
"10011111", 
"01010100", 
"10001101", 
"10010011", 
"00101110", 
"01101000", 
"01111111", 
"10010001", 
"01111111", 
"10010011", 
"10001001", 
"10001111", 
"01110010", 
"01100110", 
"11000101", 
"01111101", 
"01110111", 
"00111100", 
"10001100", 
"10101011", 
"10001110", 
"10011010", 
"10001001", 
"01110110", 
"10001110", 
"01110001", 
"01000110", 
"10010111", 
"01010100", 
"10100101", 
"01111000", 
"10011110", 
"10001001", 
"01011000", 
"11001001", 
"10011100", 
"10011001", 
"10001011", 
"10000011", 
"10011110", 
"10011101", 
"01101111", 
"01100011", 
"10000110", 
"01111011", 
"10000000", 
"01100011", 
"01111000", 
"01101110", 
"01111100", 
"10101000", 
"10001101", 
"10001100", 
"01111101", 
"10000010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_7 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_7(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
