use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_37_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_37_LAYER;

architecture Behavioral of ROM_FC_120_37_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_37: ROM_ARRAY_PESOS_FC_120 := (
"10000110", 
"10000111", 
"01100010", 
"01100111", 
"01111100", 
"01011111", 
"10000001", 
"01111001", 
"10001111", 
"01011110", 
"10011010", 
"10010111", 
"10001110", 
"10000000", 
"10010000", 
"01101111", 
"10001100", 
"01110010", 
"01011110", 
"00111101", 
"10001101", 
"10000011", 
"01100010", 
"10000010", 
"10010000", 
"10000111", 
"10000110", 
"10111101", 
"10010111", 
"01110001", 
"10000000", 
"10001010", 
"01101101", 
"01111010", 
"01110110", 
"01101100", 
"10010010", 
"01110011", 
"01001010", 
"10010010", 
"10001010", 
"01111111", 
"01101111", 
"10100001", 
"01111000", 
"01111011", 
"01101100", 
"01111001", 
"01111011", 
"11001000", 
"10000001", 
"01100010", 
"01110111", 
"01001101", 
"01110101", 
"10000110", 
"01110100", 
"01100011", 
"01110011", 
"10001100", 
"01111100", 
"01100100", 
"10010011", 
"01110001", 
"01110001", 
"01010110", 
"01111100", 
"01110100", 
"10001000", 
"01101110", 
"10001010", 
"10001100", 
"10010000", 
"10000101", 
"10001110", 
"01110000", 
"01000010", 
"10010110", 
"10000111", 
"01110001", 
"01110001", 
"01110010", 
"01111010", 
"10001010", 
"01110101", 
"10000111", 
"10010000", 
"01101101", 
"10001000", 
"01101011", 
"10001010", 
"01110111", 
"10001101", 
"01101111", 
"10000110", 
"01101111", 
"01110010", 
"10100001", 
"01100111", 
"01000100", 
"01110100", 
"01101111", 
"01011101", 
"01111001", 
"10001010", 
"01110000", 
"01110100", 
"01110111", 
"10010100", 
"10011001", 
"01110110", 
"10010011", 
"01111001", 
"01100000", 
"01101011", 
"01101111", 
"10000011", 
"10001100", 
"01111111", 
"10011010", 
"01111111", 
"01101111", 
"01111100", 
"01111111", 
"10000110", 
"10010100", 
"01111100", 
"10000100", 
"01101000", 
"01010010", 
"10001100", 
"10101101", 
"01101110", 
"01110101", 
"01110110", 
"01100101", 
"01101101", 
"01011110", 
"01110010", 
"00111001", 
"01101010", 
"01100110", 
"01111111", 
"10000010", 
"01110000", 
"10001100", 
"01100010", 
"01110110", 
"10001000", 
"10010000", 
"01111101", 
"01101111", 
"10001011", 
"10001100", 
"01110100", 
"01100101", 
"01000010", 
"01100010", 
"10000011", 
"10001000", 
"01100010", 
"10010001", 
"01111001", 
"01100100", 
"01111000", 
"10010010", 
"01011100", 
"01100110", 
"01111000", 
"01010110", 
"10010111", 
"01110001", 
"01100011", 
"10011101", 
"01110001", 
"01110101", 
"10000001", 
"10100011", 
"01010100", 
"01001110", 
"10000101", 
"10001011", 
"01111110", 
"01100011", 
"10001010", 
"01001000", 
"01111000", 
"01010111", 
"01111000", 
"10100111", 
"10001001", 
"01111110", 
"01101111", 
"10000001", 
"10000111", 
"01110111", 
"10000101", 
"01011011", 
"01110111", 
"10011001", 
"01101110", 
"10011000", 
"01110101", 
"01100100", 
"10001000", 
"01101011", 
"10000110", 
"01111111", 
"01111100", 
"10000101", 
"01110100", 
"01111101", 
"01111101", 
"01100011", 
"10000001", 
"10001101", 
"01111110", 
"10010011", 
"01101101", 
"10011000", 
"10110011", 
"01101110", 
"01111011", 
"01110001", 
"10100100", 
"10011011", 
"01011100", 
"01011101", 
"01111000", 
"01111011", 
"10000010", 
"01111001", 
"10000110", 
"01111101", 
"01101001", 
"01101110", 
"01101010", 
"10000010", 
"10001101", 
"01111011", 
"10011010", 
"01111001", 
"01111101", 
"01011001", 
"10001010", 
"10100011", 
"10010111", 
"01111011", 
"10001010", 
"01110110", 
"10000111", 
"01011001", 
"01100001", 
"01101110", 
"10001011", 
"01110111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_37: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_37(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
