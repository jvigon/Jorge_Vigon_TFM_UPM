use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_27_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_27_LAYER;

architecture Behavioral of ROM_FC_120_27_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_27: ROM_ARRAY_PESOS_FC_120 := (
"10011001", 
"01111001", 
"01101111", 
"10111110", 
"01111101", 
"01101101", 
"01001100", 
"10000100", 
"01110000", 
"10010101", 
"01100001", 
"10001011", 
"01111100", 
"10010010", 
"01110011", 
"10011001", 
"10010001", 
"01100100", 
"01110101", 
"01111100", 
"10001100", 
"01111000", 
"01011001", 
"10001011", 
"10001111", 
"10011000", 
"01111010", 
"01111101", 
"10001110", 
"01011000", 
"01110100", 
"10000011", 
"01101101", 
"01100100", 
"10000011", 
"10001011", 
"10001111", 
"10000000", 
"10001001", 
"01110100", 
"01111001", 
"10001010", 
"01110100", 
"01111111", 
"01011110", 
"10010000", 
"01110110", 
"01100001", 
"01100010", 
"01111011", 
"10101001", 
"10000010", 
"10001010", 
"10010100", 
"01110110", 
"01101111", 
"01111001", 
"01000111", 
"10000111", 
"01111100", 
"01010101", 
"01111010", 
"01110110", 
"01011111", 
"10001111", 
"01111101", 
"01110011", 
"01110100", 
"01110000", 
"01100010", 
"10010010", 
"10100110", 
"10001110", 
"10010001", 
"01011010", 
"01110001", 
"10110110", 
"10100011", 
"10001001", 
"01110111", 
"01110111", 
"01110011", 
"01101110", 
"01011001", 
"01101110", 
"10000110", 
"01110010", 
"10011101", 
"10001111", 
"01100111", 
"01111001", 
"01101001", 
"10000111", 
"10001101", 
"01111010", 
"01111000", 
"01111001", 
"01011111", 
"01111001", 
"10000001", 
"01110111", 
"01110111", 
"10000111", 
"01110001", 
"10000111", 
"10000100", 
"01101111", 
"10000001", 
"10011111", 
"10011010", 
"01101100", 
"01111011", 
"10001001", 
"01100101", 
"01111011", 
"10000011", 
"01110010", 
"10001010", 
"10001001", 
"01111100", 
"01110110", 
"10001110", 
"01111110", 
"01110010", 
"01110011", 
"10000010", 
"01110110", 
"10001000", 
"10001111", 
"01101110", 
"10010100", 
"01101010", 
"01111111", 
"01101110", 
"10101001", 
"10010010", 
"10001011", 
"01110011", 
"10101101", 
"10000111", 
"11011110", 
"01001100", 
"10000110", 
"01110011", 
"10010101", 
"10101111", 
"10000010", 
"00110111", 
"01111011", 
"01111000", 
"10001100", 
"01110011", 
"10001101", 
"01111001", 
"01111001", 
"01110100", 
"10010010", 
"01111101", 
"01101110", 
"10000100", 
"01110101", 
"10100011", 
"01111000", 
"01001101", 
"01101111", 
"01111010", 
"01111010", 
"01101001", 
"10010011", 
"10011000", 
"10000011", 
"01100101", 
"01110000", 
"01110011", 
"10000010", 
"10000101", 
"01101100", 
"01100101", 
"01101000", 
"11000011", 
"01111100", 
"01110000", 
"10000001", 
"10000100", 
"01111000", 
"10000110", 
"01110001", 
"10001001", 
"01110011", 
"10100000", 
"10001010", 
"01110011", 
"01111001", 
"10000110", 
"10010000", 
"10110110", 
"01110111", 
"10001111", 
"01111101", 
"10011111", 
"01110000", 
"10100111", 
"10100010", 
"01001110", 
"10001000", 
"01010001", 
"01110010", 
"10001101", 
"10001001", 
"10010000", 
"10000000", 
"01101100", 
"10001100", 
"10000100", 
"01110010", 
"10011110", 
"01101111", 
"10000010", 
"10000001", 
"01101011", 
"01101110", 
"01101100", 
"10000101", 
"10001000", 
"01101110", 
"10000100", 
"10000100", 
"01011010", 
"01110111", 
"01100011", 
"01100000", 
"10010010", 
"10000010", 
"01101110", 
"01100101", 
"10100010", 
"01100000", 
"01101011", 
"10001100", 
"01111101", 
"01101100", 
"01110011", 
"01111010", 
"10011001", 
"01101101", 
"01111000", 
"10010111", 
"01110110", 
"10001101", 
"10000101", 
"01100010", 
"10001111", 
"01010101", 
"10001101", 
"10000010", 
"01110010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_27: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_27(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
