use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_11_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_11_LAYER;

architecture Behavioral of ROM_FC_120_11_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_11: ROM_ARRAY_PESOS_FC_120 := (
"01110111", 
"01101010", 
"10000110", 
"01100001", 
"01011011", 
"01010010", 
"10001000", 
"10011000", 
"01111001", 
"01110100", 
"01011110", 
"10000100", 
"10011011", 
"01101100", 
"01100000", 
"10010111", 
"00111001", 
"01100100", 
"10001000", 
"01010100", 
"10101001", 
"00010010", 
"10001101", 
"01101100", 
"10001101", 
"01110001", 
"10010001", 
"01101111", 
"10001101", 
"01001101", 
"01111000", 
"10000111", 
"00110110", 
"10001101", 
"10100001", 
"01010101", 
"10001011", 
"00100100", 
"01101110", 
"00101101", 
"01110001", 
"10010011", 
"10000110", 
"01111100", 
"10010001", 
"01100110", 
"10011011", 
"10001010", 
"00111000", 
"10010011", 
"01101111", 
"01100100", 
"10010101", 
"10001100", 
"00100111", 
"00110101", 
"01111110", 
"10011100", 
"10000010", 
"10011000", 
"01100000", 
"10010010", 
"10001000", 
"10000010", 
"10001011", 
"10001101", 
"10100111", 
"01110001", 
"10000110", 
"10100101", 
"10001000", 
"01101010", 
"01111001", 
"01111100", 
"10001110", 
"01001100", 
"01100101", 
"01001000", 
"01111110", 
"01101100", 
"10011110", 
"01111111", 
"01111000", 
"01110010", 
"01100010", 
"10001001", 
"10001011", 
"01100111", 
"10000000", 
"01111001", 
"01011110", 
"10010001", 
"01011000", 
"01111011", 
"10001010", 
"10000000", 
"01100100", 
"10100101", 
"10000100", 
"01101011", 
"01111111", 
"01110110", 
"01101001", 
"01011011", 
"01011100", 
"01010101", 
"01101010", 
"10001000", 
"01001000", 
"10010101", 
"01111011", 
"01101011", 
"10001111", 
"11001010", 
"01011100", 
"01001000", 
"01110111", 
"01111111", 
"11001111", 
"01100001", 
"10000000", 
"01000010", 
"10100000", 
"10101011", 
"01111111", 
"01011001", 
"01111101", 
"10000111", 
"10000100", 
"10001101", 
"01111101", 
"10011100", 
"01101111", 
"10011111", 
"01101110", 
"10111100", 
"01111100", 
"10001100", 
"10001111", 
"01101001", 
"00111111", 
"01110000", 
"01101010", 
"10000011", 
"10100000", 
"01101001", 
"10001001", 
"10100100", 
"01110001", 
"01111010", 
"10000111", 
"10100101", 
"10000110", 
"01101001", 
"01101010", 
"01101011", 
"01100001", 
"10010011", 
"01101011", 
"01101101", 
"10011011", 
"01011101", 
"10001011", 
"01000100", 
"10000001", 
"01111111", 
"10010100", 
"10100101", 
"01110001", 
"10000100", 
"10001000", 
"10010111", 
"01101111", 
"01010010", 
"10100000", 
"10010111", 
"10011000", 
"01101110", 
"01010100", 
"00100101", 
"10001010", 
"01110110", 
"01100010", 
"10010111", 
"10010000", 
"01111010", 
"10000101", 
"10001001", 
"01100011", 
"00111101", 
"10001000", 
"10000101", 
"01101010", 
"01011000", 
"01101110", 
"10001100", 
"01101101", 
"01110100", 
"10001000", 
"10100000", 
"01101011", 
"01101101", 
"01111011", 
"10100001", 
"01111000", 
"01110011", 
"10001010", 
"01111000", 
"11001111", 
"00111101", 
"01011111", 
"10001100", 
"01100101", 
"01110000", 
"10011110", 
"01111010", 
"10100000", 
"10000011", 
"01101110", 
"10001110", 
"01010011", 
"10101110", 
"01111100", 
"01011000", 
"10100111", 
"01010000", 
"01011101", 
"01011111", 
"01101001", 
"01011011", 
"01101101", 
"10100010", 
"10010111", 
"10001111", 
"01100010", 
"01100101", 
"10000010", 
"01001011", 
"10001111", 
"01111001", 
"01101100", 
"00110101", 
"01111110", 
"01000011", 
"10010001", 
"01101110", 
"01001100", 
"10100011", 
"10001100", 
"10000001", 
"01000110", 
"01011110", 
"01111011", 
"01010110", 
"10001001", 
"01111011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_11: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_11(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
