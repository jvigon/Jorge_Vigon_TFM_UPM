use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_109_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_109_LAYER;

architecture Behavioral of ROM_FC_120_109_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_109: ROM_ARRAY_PESOS_FC_120 := (
"01110001", 
"10001101", 
"01101000", 
"10001100", 
"11000000", 
"01100000", 
"01111010", 
"00111100", 
"10001001", 
"10100100", 
"01101100", 
"10100100", 
"01111111", 
"01100010", 
"01110001", 
"01111101", 
"10001001", 
"01011010", 
"01011010", 
"01111011", 
"01100110", 
"11011100", 
"01110101", 
"10001100", 
"10111100", 
"01011110", 
"10011010", 
"01100100", 
"00101111", 
"10001010", 
"01111000", 
"01110111", 
"10000010", 
"01000000", 
"01111010", 
"10011001", 
"10011010", 
"01110011", 
"01011111", 
"10101000", 
"10000001", 
"01111100", 
"01011000", 
"01101110", 
"01011001", 
"10100000", 
"10000110", 
"10010001", 
"01101010", 
"01001101", 
"00111001", 
"10000010", 
"01111010", 
"10110010", 
"01110110", 
"01100001", 
"10001100", 
"00111001", 
"01001100", 
"01111100", 
"01000001", 
"01010101", 
"01101111", 
"10001001", 
"10000011", 
"01011100", 
"01011110", 
"10001100", 
"01100000", 
"10010001", 
"01100011", 
"01100110", 
"10010011", 
"10000111", 
"01101001", 
"01110000", 
"01101010", 
"01011111", 
"01111100", 
"01111011", 
"01101111", 
"00110001", 
"01001011", 
"01110111", 
"10000010", 
"11010001", 
"01101011", 
"01010100", 
"10101111", 
"01010111", 
"01110101", 
"10010100", 
"01100110", 
"10001001", 
"10000001", 
"01111001", 
"10101101", 
"01101111", 
"10000101", 
"01101110", 
"01110110", 
"01111111", 
"01010010", 
"01101101", 
"10100101", 
"01111100", 
"01100100", 
"01100010", 
"01010011", 
"11100100", 
"01110101", 
"10000001", 
"10001110", 
"01110001", 
"01000010", 
"00111101", 
"01110001", 
"10010000", 
"10010111", 
"01100111", 
"01111011", 
"00100010", 
"01011010", 
"10110011", 
"01111000", 
"10100111", 
"01110001", 
"10001010", 
"01111011", 
"01000000", 
"01111001", 
"01110001", 
"01101111", 
"10010111", 
"01110100", 
"01110010", 
"01111111", 
"01100011", 
"10001111", 
"01111111", 
"01101110", 
"10111000", 
"01111000", 
"01111101", 
"10010100", 
"01010000", 
"01011010", 
"10010111", 
"01111001", 
"10011100", 
"01001100", 
"10001001", 
"10100101", 
"01001101", 
"01001001", 
"01000100", 
"01100011", 
"10110111", 
"01111000", 
"10001110", 
"01100110", 
"01100101", 
"10001010", 
"10010100", 
"01111000", 
"10011000", 
"01010100", 
"01111110", 
"10110100", 
"01101100", 
"10001100", 
"01101100", 
"10001100", 
"11001110", 
"01111011", 
"10001001", 
"10001000", 
"01001001", 
"10011000", 
"01110101", 
"10010010", 
"01010011", 
"01111000", 
"01001101", 
"01101001", 
"01100001", 
"01000010", 
"01110101", 
"10110101", 
"10010101", 
"10000110", 
"10010011", 
"01111100", 
"10100010", 
"00111101", 
"01111001", 
"01101001", 
"11011011", 
"11000001", 
"10100001", 
"10001110", 
"01101100", 
"10010110", 
"01110111", 
"00101011", 
"01111010", 
"01101101", 
"01111011", 
"10001000", 
"10100000", 
"01110110", 
"01011001", 
"10001001", 
"10000100", 
"01011111", 
"01011010", 
"01110101", 
"01011101", 
"00111111", 
"01110011", 
"01011001", 
"01111010", 
"01101011", 
"10000101", 
"01010011", 
"01111110", 
"00110101", 
"01100100", 
"10000111", 
"01110100", 
"01111010", 
"01010011", 
"10000000", 
"01100100", 
"01111000", 
"01111001", 
"01100000", 
"01010111", 
"01111100", 
"10001010", 
"01011100", 
"01111101", 
"01101110", 
"10001110", 
"01111100", 
"01011111", 
"10011011", 
"01100001", 
"01111101", 
"01111010", 
"01100001", 
"10001101", 
"10000110", 
"11000000", 
"10001111", 
"01110110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_109 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_109(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
