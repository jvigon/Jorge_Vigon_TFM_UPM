use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_78_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_78_LAYER;

architecture Behavioral of ROM_FC_84_78_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_78: ROM_ARRAY_PESOS_FC_84 := (
"01101011", 
"10000001", 
"10000010", 
"01011001", 
"01110101", 
"10010110", 
"01101111", 
"10011100", 
"01100101", 
"10010110", 
"10100100", 
"01010010", 
"01101010", 
"01110100", 
"01101001", 
"10100110", 
"10000000", 
"01101000", 
"10011011", 
"10100100", 
"01110111", 
"10011001", 
"10000000", 
"01111000", 
"10001101", 
"01011011", 
"01110001", 
"10010010", 
"10110010", 
"10010100", 
"01111100", 
"10001010", 
"01100110", 
"11001100", 
"01110110", 
"00111111", 
"01111000", 
"01110101", 
"10100110", 
"01101111", 
"01011010", 
"10010101", 
"00011010", 
"10000000", 
"10000110", 
"01111111", 
"01101110", 
"01110100", 
"00111001", 
"10011001", 
"01100111", 
"10101001", 
"10010101", 
"01001100", 
"10100001", 
"10111100", 
"10010111", 
"01111000", 
"01100111", 
"10100101", 
"10010010", 
"01111001", 
"01100001", 
"01010000", 
"01111001", 
"01101101", 
"10010001", 
"01011001", 
"10010101", 
"10001010", 
"01011111", 
"01100000", 
"01011111", 
"01110001", 
"01111101", 
"01110010", 
"01100010", 
"10100111", 
"01111000", 
"10000101", 
"01101110", 
"01101110", 
"10011000", 
"10101001", 
"01101100", 
"01100001", 
"10011000", 
"01101010", 
"01111100", 
"11000110", 
"01011110", 
"11010001", 
"01111011", 
"10000100", 
"01111100", 
"01101111", 
"10000001", 
"10000110", 
"01011010", 
"01110001", 
"10000111", 
"10101011", 
"01101111", 
"01110000", 
"00110011", 
"10100010", 
"10000010", 
"01111101", 
"10000101", 
"11011000", 
"01101101", 
"10101011", 
"01110110", 
"01001101", 
"10000000", 
"10011000", 
"10100110", 
"01001001", 
"10001011", 
"10101000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_78: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_78(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
