use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_36_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_36_LAYER;

architecture Behavioral of ROM_FC_120_36_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_36: ROM_ARRAY_PESOS_FC_120 := (
"01101111", 
"10100100", 
"01100000", 
"00101010", 
"10001001", 
"01111111", 
"00101010", 
"01101011", 
"01101011", 
"10011010", 
"01011101", 
"11111111", 
"10000010", 
"01110110", 
"10000101", 
"01111111", 
"10000100", 
"10101110", 
"01010011", 
"01111010", 
"01011010", 
"10101000", 
"01001110", 
"01100101", 
"10000101", 
"01010000", 
"01100110", 
"10111101", 
"01101101", 
"01111001", 
"10010100", 
"01101111", 
"10001001", 
"01111101", 
"01000011", 
"10010111", 
"10000010", 
"01011100", 
"10000100", 
"10001011", 
"10000010", 
"01000101", 
"10001010", 
"01100111", 
"01010111", 
"10011000", 
"01111000", 
"01110110", 
"01110001", 
"01010000", 
"10010001", 
"10010111", 
"10001011", 
"01011101", 
"10001001", 
"10101010", 
"01111100", 
"01011111", 
"01101000", 
"01000011", 
"00111110", 
"01101010", 
"10001100", 
"01111100", 
"01100100", 
"00100100", 
"01010110", 
"01100000", 
"10000111", 
"00110100", 
"00100101", 
"10000000", 
"01101101", 
"01111100", 
"01101011", 
"10010001", 
"10010011", 
"10111010", 
"01101101", 
"10000000", 
"01101001", 
"01111011", 
"00111010", 
"01001000", 
"10000111", 
"01000000", 
"01011101", 
"01110001", 
"10000010", 
"10101011", 
"01011100", 
"01011011", 
"01111001", 
"01100111", 
"01110000", 
"01111101", 
"10001111", 
"01110001", 
"01111010", 
"01111100", 
"01101101", 
"01011110", 
"01100111", 
"10010110", 
"01111001", 
"01111110", 
"01111000", 
"01100111", 
"00110111", 
"01010010", 
"10000100", 
"10000010", 
"01011100", 
"01001110", 
"01110000", 
"01101101", 
"01111111", 
"01000110", 
"01100110", 
"01100011", 
"10001100", 
"01101010", 
"01101110", 
"01110111", 
"01001000", 
"01110111", 
"10001100", 
"10000101", 
"01110000", 
"01010000", 
"01001100", 
"00101111", 
"01101100", 
"01110001", 
"01011100", 
"10000111", 
"01101110", 
"10110011", 
"01101100", 
"01110000", 
"10010111", 
"01010110", 
"01111011", 
"01101001", 
"01110110", 
"10010001", 
"00110101", 
"00101111", 
"10000101", 
"01011001", 
"10001100", 
"10110010", 
"01111001", 
"10001001", 
"00010110", 
"10001011", 
"10011011", 
"01101011", 
"10000000", 
"01101110", 
"01111110", 
"10100001", 
"01010111", 
"01000010", 
"10001011", 
"10010101", 
"01111010", 
"10010011", 
"01100011", 
"01011100", 
"00111101", 
"10001110", 
"01011011", 
"10010011", 
"01111000", 
"01111011", 
"10011010", 
"10011001", 
"01011011", 
"01000100", 
"10001001", 
"01111010", 
"10100000", 
"01001111", 
"01111000", 
"10100100", 
"01101000", 
"01101001", 
"10000011", 
"01111000", 
"10000111", 
"01111000", 
"01100110", 
"01010100", 
"10001111", 
"01000010", 
"10000001", 
"10001100", 
"01111110", 
"01101111", 
"10000011", 
"10000011", 
"01101011", 
"10000000", 
"01001100", 
"01101011", 
"01110010", 
"01111001", 
"01010101", 
"10111001", 
"01111001", 
"10000001", 
"10001000", 
"01010010", 
"01101010", 
"01110100", 
"10001110", 
"01111100", 
"10010000", 
"01111110", 
"01100001", 
"01111101", 
"01110000", 
"01110100", 
"10100011", 
"10001010", 
"01111001", 
"01010001", 
"10000000", 
"01111011", 
"01100001", 
"01111010", 
"01100001", 
"01111111", 
"01001001", 
"01001000", 
"10100111", 
"01101101", 
"01111111", 
"01110100", 
"10001110", 
"01110101", 
"01101100", 
"01101011", 
"01101111", 
"01111111", 
"01100101", 
"01110110", 
"10001100", 
"01111001", 
"10001011", 
"01101111", 
"01101000", 
"01111101", 
"01110111", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_36: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_36(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
