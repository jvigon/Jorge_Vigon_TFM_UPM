use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_13_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_13_LAYER;

architecture Behavioral of ROM_FC_84_13_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_13: ROM_ARRAY_PESOS_FC_84 := (
"00110011", 
"01111011", 
"10001101", 
"10000110", 
"10010010", 
"10000110", 
"01100111", 
"01011001", 
"01110110", 
"01010011", 
"10110000", 
"01101000", 
"01011001", 
"01110010", 
"01101001", 
"10001110", 
"10000010", 
"01110111", 
"01001100", 
"01011011", 
"01100100", 
"10111010", 
"01110000", 
"10011110", 
"01101001", 
"01111010", 
"10001110", 
"01101000", 
"10000101", 
"10010010", 
"01111001", 
"01000101", 
"01100101", 
"10000101", 
"01100101", 
"01001000", 
"10101001", 
"10010011", 
"10101001", 
"01010010", 
"01110110", 
"00110101", 
"01010011", 
"10001101", 
"01100001", 
"01011001", 
"10010101", 
"01101010", 
"01100000", 
"10001010", 
"01111110", 
"01110010", 
"01110111", 
"01100011", 
"10001000", 
"01101010", 
"10000001", 
"01110111", 
"00111101", 
"10100000", 
"10000011", 
"01011100", 
"01101100", 
"01011010", 
"10001011", 
"10110001", 
"01010010", 
"01110000", 
"10001111", 
"10011111", 
"10100010", 
"00110001", 
"01110011", 
"01001101", 
"01111000", 
"10010010", 
"10001110", 
"01101100", 
"01111011", 
"01111101", 
"01110100", 
"10001001", 
"10010001", 
"01110110", 
"01111110", 
"01100111", 
"01110111", 
"10000100", 
"10010000", 
"10001011", 
"10010001", 
"10100001", 
"10011000", 
"01101110", 
"01100011", 
"01001110", 
"01101001", 
"10001000", 
"10010111", 
"01110010", 
"10010110", 
"10100001", 
"01111111", 
"10001111", 
"00111011", 
"01110010", 
"10010001", 
"10000110", 
"01110011", 
"11001001", 
"01100010", 
"10001001", 
"10010101", 
"10000001", 
"01111101", 
"01110111", 
"10010100", 
"01000111", 
"10001010", 
"01100011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_13 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_13(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
