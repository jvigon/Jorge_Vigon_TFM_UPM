use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_4_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_4_LAYER;

architecture Behavioral of ROM_FC_120_4_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_4: ROM_ARRAY_PESOS_FC_120 := (
"01111111", 
"01000011", 
"10101111", 
"10011100", 
"10001111", 
"01101110", 
"01001101", 
"01100010", 
"01110110", 
"10000110", 
"10011001", 
"01011100", 
"10010110", 
"01110101", 
"01110101", 
"10110110", 
"01100111", 
"00111111", 
"01100110", 
"10110001", 
"01111011", 
"01101001", 
"10101111", 
"01100100", 
"10001101", 
"01001010", 
"01100100", 
"01100011", 
"01101111", 
"01110011", 
"01110100", 
"10001001", 
"10001101", 
"01111000", 
"01111011", 
"01111111", 
"01101011", 
"10001100", 
"01010001", 
"01011111", 
"10001100", 
"10010100", 
"10000001", 
"01001111", 
"10010111", 
"01100100", 
"10001001", 
"10010001", 
"10001010", 
"00111010", 
"10000100", 
"10100010", 
"01101011", 
"01000000", 
"10001010", 
"01101111", 
"01101111", 
"10001101", 
"01101011", 
"00010001", 
"10110000", 
"01101000", 
"10000011", 
"10011000", 
"01110011", 
"01111010", 
"10000101", 
"10011101", 
"01101100", 
"10101100", 
"01011100", 
"01110100", 
"10000100", 
"10000101", 
"10100111", 
"10011100", 
"01001111", 
"01101111", 
"01111001", 
"10000000", 
"01101110", 
"01111111", 
"01101000", 
"01010110", 
"10001011", 
"01100001", 
"01101100", 
"01100010", 
"10000010", 
"10000010", 
"01000010", 
"10011001", 
"01101011", 
"01111110", 
"10000010", 
"10001011", 
"01100101", 
"10010000", 
"10000010", 
"01111011", 
"10000101", 
"01111001", 
"01011001", 
"01001001", 
"01111100", 
"10001111", 
"01101010", 
"01111011", 
"01110111", 
"01011001", 
"01100111", 
"01111000", 
"01000111", 
"01111011", 
"01101010", 
"01100010", 
"10010010", 
"01000101", 
"01010101", 
"01010000", 
"01111101", 
"01101010", 
"01101101", 
"01101110", 
"10001101", 
"01010101", 
"10000011", 
"10001100", 
"10000000", 
"01101100", 
"01110011", 
"10101111", 
"01101011", 
"10110011", 
"01111100", 
"10001011", 
"10000100", 
"10000101", 
"01101100", 
"01100110", 
"01111101", 
"10000100", 
"01111001", 
"01111011", 
"01100100", 
"01110110", 
"01100011", 
"10101000", 
"01111110", 
"10000011", 
"10010101", 
"10010100", 
"10000101", 
"01010000", 
"01100010", 
"01011010", 
"10000001", 
"10001001", 
"10000110", 
"01110001", 
"01100001", 
"01010110", 
"01010100", 
"01000100", 
"01101001", 
"01101000", 
"10001010", 
"01110011", 
"01101111", 
"01100011", 
"01111101", 
"10000010", 
"10010011", 
"01111001", 
"10000000", 
"01111101", 
"01100001", 
"01101110", 
"10000100", 
"00110001", 
"01101000", 
"01000110", 
"10101011", 
"01011001", 
"10000110", 
"10001011", 
"01100111", 
"01011001", 
"10010001", 
"01111111", 
"10001011", 
"01111001", 
"01111100", 
"10001110", 
"01010111", 
"01100000", 
"01101000", 
"01100110", 
"01100001", 
"01100100", 
"01101101", 
"01100001", 
"01101001", 
"10011111", 
"01111001", 
"01100110", 
"10001001", 
"10001000", 
"01101101", 
"10000011", 
"01101101", 
"01110011", 
"01110110", 
"10000100", 
"01101000", 
"01011001", 
"01101100", 
"01111010", 
"01101110", 
"01010011", 
"01100110", 
"10100001", 
"10001001", 
"01111110", 
"01110100", 
"01100101", 
"10001110", 
"10000110", 
"01101111", 
"01101111", 
"10001111", 
"01101101", 
"01110111", 
"01110101", 
"01110010", 
"01001110", 
"10101101", 
"01011001", 
"10000111", 
"10000011", 
"01100010", 
"01001011", 
"01111001", 
"10100011", 
"10000111", 
"01101100", 
"01011000", 
"01011101", 
"10000011", 
"01111100", 
"01100001", 
"01011101", 
"10011000", 
"01110101", 
"01110100", 
"01111011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_4 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_4(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
