use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_18_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_18_LAYER;

architecture Behavioral of ROM_FC_84_18_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_18: ROM_ARRAY_PESOS_FC_84 := (
"01110100", 
"01001110", 
"01110001", 
"10001000", 
"10110101", 
"01111011", 
"01111011", 
"10101110", 
"10000110", 
"01110011", 
"01110010", 
"10100001", 
"01010110", 
"10111010", 
"10011010", 
"10001011", 
"01010101", 
"10001011", 
"10100000", 
"01110000", 
"10101100", 
"10001010", 
"01011111", 
"01100111", 
"01101000", 
"10100110", 
"10001011", 
"01000110", 
"01100011", 
"01011111", 
"10001011", 
"10101100", 
"10000000", 
"10001101", 
"01110011", 
"10000101", 
"01100100", 
"01101000", 
"10100110", 
"10000001", 
"01100110", 
"10000001", 
"10110010", 
"01000110", 
"00100101", 
"01101010", 
"01110101", 
"10001000", 
"01001000", 
"10001110", 
"01101101", 
"01101110", 
"01111011", 
"01001011", 
"01110101", 
"01110111", 
"10011000", 
"10100000", 
"10100000", 
"01010100", 
"01110010", 
"01110011", 
"01100011", 
"10000110", 
"01111111", 
"01000111", 
"01010001", 
"10010001", 
"01110100", 
"00111100", 
"01111101", 
"10000110", 
"00111011", 
"01100000", 
"10010100", 
"01111000", 
"10110001", 
"01100100", 
"01110001", 
"01110110", 
"10000010", 
"01110011", 
"01010011", 
"01110111", 
"10000110", 
"10000010", 
"01101010", 
"10100011", 
"10000100", 
"10101011", 
"10001111", 
"10101000", 
"10001001", 
"01101010", 
"01111110", 
"10011101", 
"10001110", 
"10010011", 
"10001001", 
"01101000", 
"01110001", 
"01110111", 
"10001011", 
"01100111", 
"01010101", 
"01100101", 
"10000010", 
"01101011", 
"10000111", 
"00110111", 
"10110010", 
"01100000", 
"10000111", 
"01000111", 
"01100001", 
"10110010", 
"01100101", 
"01011001", 
"10000011", 
"01100011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_18 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_18(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
