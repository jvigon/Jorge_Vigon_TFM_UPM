use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity ROM_FC_120_0_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_0_LAYER;

architecture Behavioral of ROM_FC_120_0_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120_0 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
-- Directiva para forzar el uso de Block RAM

--CONSTANT ROM_FC_120_0: ROM_ARRAY_PESOS_FC_120_0 := (
signal ROM_FC_120_0: ROM_ARRAY_PESOS_FC_120_0 := (
"10011010", 
"10011010", 
"01010100", 
"01010100", 
"01100111", 
"10110000", 
"10100011", 
"10010110", 
"10000111", 
"01010000", 
"01011111", 
"10110001", 
"00101111", 
"10111000", 
"01111001", 
"01110011", 
"10001110", 
"01110111", 
"01110100", 
"01011001", 
"01101001", 
"10100110", 
"10010010", 
"01111100", 
"01111010", 
"01101011", 
"01101000", 
"10000100", 
"01010010", 
"10110101", 
"01110110", 
"10001000", 
"01110101", 
"10111100", 
"10000011", 
"01110110", 
"10010000", 
"10010000", 
"10001110", 
"01011111", 
"10000010", 
"01001010", 
"10010101", 
"10001111", 
"01110010", 
"01111110", 
"10001110", 
"01111000", 
"10010000", 
"01101101", 
"01100100", 
"10000101", 
"10000110", 
"10110101", 
"01111011", 
"10000100", 
"10010000", 
"01010010", 
"01111111", 
"01110100", 
"01000110", 
"10000101", 
"01101101", 
"10001110", 
"01111010", 
"01110100", 
"10000010", 
"01110100", 
"10101000", 
"10101101", 
"10111100", 
"10010101", 
"10001011", 
"01000100", 
"01111110", 
"01010111", 
"11001110", 
"01010101", 
"10010100", 
"01110101", 
"10101000", 
"10000010", 
"10001010", 
"01100100", 
"10010100", 
"10011001", 
"10010100", 
"10100001", 
"01111011", 
"01111101", 
"10010000", 
"01110011", 
"10000001", 
"01001110", 
"01110101", 
"10001100", 
"01010111", 
"01111001", 
"10011111", 
"10001110", 
"01110111", 
"01100010", 
"10101011", 
"10001110", 
"01111110", 
"01010000", 
"01111110", 
"10101011", 
"01101110", 
"01100101", 
"01110111", 
"01110101", 
"10100101", 
"01000011", 
"10001001", 
"10100100", 
"10010010", 
"10011101", 
"10001011", 
"01111111", 
"10001001", 
"01101010", 
"10010110", 
"01101110", 
"01101101", 
"10001110", 
"01110110", 
"10001101", 
"01100000", 
"01011011", 
"10001000", 
"10000101", 
"10000010", 
"01010010", 
"10101001", 
"01110110", 
"10001000", 
"10011000", 
"10101011", 
"01001110", 
"01110111", 
"01011010", 
"10000111", 
"10000101", 
"10001100", 
"01111100", 
"10100001", 
"10010110", 
"01110000", 
"01001101", 
"01101100", 
"10001111", 
"10000111", 
"01101000", 
"10100010", 
"01111010", 
"10100100", 
"01110011", 
"10001110", 
"10001011", 
"10000011", 
"01111010", 
"10011111", 
"10100001", 
"10001111", 
"01010010", 
"10100000", 
"01010111", 
"10010001", 
"01101010", 
"01011110", 
"10010000", 
"01110111", 
"10010111", 
"10010011", 
"10000111", 
"01110011", 
"01011000", 
"10010011", 
"10100011", 
"01111110", 
"10100000", 
"10010001", 
"10001000", 
"10010101", 
"10010011", 
"10001010", 
"01111100", 
"01110111", 
"01010111", 
"01111011", 
"01110101", 
"01111100", 
"10000100", 
"01100001", 
"01110101", 
"10001100", 
"10000010", 
"10001110", 
"01110110", 
"01110100", 
"10010111", 
"01110001", 
"10010000", 
"01100110", 
"10100101", 
"10001110", 
"10001010", 
"01111011", 
"10100001", 
"10010011", 
"01110100", 
"10000011", 
"01011110", 
"01011000", 
"01000000", 
"10000101", 
"10010011", 
"10001110", 
"10011101", 
"00111110", 
"01111100", 
"01110010", 
"10010010", 
"10000000", 
"10011111", 
"01111100", 
"01111100", 
"01101101", 
"01101111", 
"01001011", 
"01010001", 
"10010000", 
"10010101", 
"10001001", 
"01111001", 
"01111010", 
"01111000", 
"10010101", 
"01110101", 
"01011110", 
"10000001", 
"10000110", 
"01101100", 
"10001010", 
"01111110", 
"01001111", 
"01011000", 
"10001001", 
"10110101", 
"10100000", 
"01100000", 
"10010111", 
"10000110", 
"10001001", 
"10000110"
);
 
attribute rom_style : string;
attribute rom_style of ROM_FC_120_0 : signal is "block";
begin 


process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_0(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
