use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_62_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_62_LAYER;

architecture Behavioral of ROM_FC_120_62_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_62: ROM_ARRAY_PESOS_FC_120 := (
"01011110", 
"01101000", 
"01110011", 
"10011000", 
"01111101", 
"01101001", 
"01001111", 
"01100100", 
"10000000", 
"01111010", 
"10000111", 
"01100100", 
"01110000", 
"10011000", 
"10010110", 
"01110011", 
"01111000", 
"01011010", 
"01100011", 
"01110110", 
"01101001", 
"01110100", 
"01101101", 
"01101111", 
"10000010", 
"01110101", 
"01001111", 
"01101100", 
"01011110", 
"10001000", 
"01101010", 
"10001110", 
"01010010", 
"01110010", 
"01111011", 
"01110011", 
"10001001", 
"01111010", 
"10000010", 
"01110011", 
"10000111", 
"01110000", 
"01011010", 
"01101110", 
"01111100", 
"01011100", 
"10000011", 
"10001100", 
"01101000", 
"01111111", 
"01110011", 
"01011110", 
"10000111", 
"01100110", 
"10001101", 
"01110011", 
"01110010", 
"01111001", 
"10001110", 
"10001000", 
"01011110", 
"01100110", 
"10011111", 
"01110110", 
"01011101", 
"01110000", 
"10010001", 
"10100101", 
"01101101", 
"10000000", 
"01111000", 
"01011111", 
"01111110", 
"01010101", 
"10000000", 
"10010011", 
"10001010", 
"10000010", 
"01011010", 
"10000010", 
"01011000", 
"01011111", 
"01111011", 
"01111101", 
"01100101", 
"01101000", 
"01011100", 
"01110010", 
"01110011", 
"01101110", 
"01110110", 
"01111110", 
"01110110", 
"01111100", 
"10000100", 
"10010001", 
"01111010", 
"01101011", 
"01111010", 
"01110001", 
"01011101", 
"01110001", 
"10000011", 
"01101101", 
"01111111", 
"10001000", 
"01010000", 
"01110000", 
"10000101", 
"01111011", 
"10000011", 
"10001001", 
"01101000", 
"01001111", 
"10001000", 
"01111010", 
"01110010", 
"01110001", 
"01111100", 
"10001000", 
"01101100", 
"01100100", 
"10001001", 
"01111000", 
"01110010", 
"01011101", 
"01110110", 
"10001000", 
"01001011", 
"10000011", 
"01100011", 
"10011110", 
"01100110", 
"01111011", 
"01110001", 
"01111000", 
"10011011", 
"01100010", 
"10011101", 
"01011111", 
"01110010", 
"10000010", 
"10001010", 
"10010000", 
"01110100", 
"10000010", 
"10010000", 
"01111000", 
"01100100", 
"01100010", 
"01111000", 
"01011011", 
"01110100", 
"10000111", 
"01110001", 
"01101100", 
"01101001", 
"01110000", 
"01110011", 
"01110000", 
"01100110", 
"10010011", 
"01101010", 
"10001100", 
"01111000", 
"01110011", 
"10000111", 
"10001001", 
"01111100", 
"01110001", 
"01100001", 
"01111000", 
"01111001", 
"01100110", 
"01110010", 
"01111000", 
"01110001", 
"01101001", 
"01100001", 
"01101001", 
"10001001", 
"01101001", 
"10010011", 
"01011100", 
"01110011", 
"01010101", 
"10001001", 
"10000101", 
"01101000", 
"01010110", 
"01111001", 
"01110101", 
"01111001", 
"01111001", 
"01111101", 
"01111010", 
"01110110", 
"01111101", 
"01111001", 
"01101111", 
"10001000", 
"01001111", 
"10001110", 
"01111111", 
"01100111", 
"01100101", 
"01111001", 
"01111100", 
"01101100", 
"01011011", 
"01101110", 
"10000000", 
"10000001", 
"01101011", 
"01111001", 
"01111100", 
"10000010", 
"01110100", 
"01101001", 
"01111111", 
"01111101", 
"01001001", 
"10001101", 
"10000110", 
"01110011", 
"01110100", 
"10000010", 
"01101100", 
"01110010", 
"01110000", 
"01101100", 
"01100110", 
"10000010", 
"01100010", 
"01100110", 
"01100100", 
"10000110", 
"10001101", 
"10000011", 
"10001110", 
"10001111", 
"01111010", 
"01111101", 
"01111011", 
"01110001", 
"01101001", 
"01111001", 
"10001100", 
"01110100", 
"01110000", 
"01110011", 
"01110101", 
"01110101", 
"01111001", 
"10001101", 
"10001111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_62: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_62(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
