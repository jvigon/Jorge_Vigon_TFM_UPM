use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_21_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_21_LAYER;

architecture Behavioral of ROM_FC_120_21_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_21: ROM_ARRAY_PESOS_FC_120 := (
"10000100", 
"01110010", 
"01101100", 
"01000111", 
"01100001", 
"10001001", 
"01101011", 
"01110001", 
"01110111", 
"00011001", 
"01100110", 
"01100000", 
"01101100", 
"01100100", 
"01111110", 
"10001011", 
"01111100", 
"01100100", 
"01001100", 
"01111001", 
"01101000", 
"10100011", 
"10000110", 
"10001010", 
"10000011", 
"00111100", 
"10100010", 
"01001000", 
"01001101", 
"01010110", 
"10001101", 
"10000111", 
"10010010", 
"01000011", 
"00111011", 
"10000001", 
"01110111", 
"10100111", 
"01111110", 
"10101111", 
"01111100", 
"10100110", 
"10011100", 
"10110001", 
"01101011", 
"10110011", 
"01110100", 
"10001011", 
"01111000", 
"01100000", 
"01100000", 
"01101001", 
"01101100", 
"10001111", 
"10011011", 
"10111110", 
"10000011", 
"10011101", 
"01001111", 
"10101010", 
"01100001", 
"01111101", 
"01111110", 
"10011111", 
"01111110", 
"10011001", 
"00110000", 
"01111110", 
"10000100", 
"10000010", 
"10000101", 
"01110110", 
"10001111", 
"01100100", 
"01010011", 
"01011011", 
"01101000", 
"01101101", 
"01111001", 
"01100110", 
"01101100", 
"10000111", 
"00111010", 
"00100100", 
"10000000", 
"01111101", 
"10101101", 
"10000110", 
"01110110", 
"01110110", 
"01011110", 
"00111110", 
"01110111", 
"01011011", 
"01110100", 
"01101111", 
"01110011", 
"10001101", 
"01010111", 
"01010110", 
"01111000", 
"01111001", 
"01110100", 
"01101100", 
"01110011", 
"10110100", 
"10101000", 
"01000101", 
"11000010", 
"01100000", 
"01111111", 
"01101100", 
"10000101", 
"01010100", 
"01011010", 
"00110010", 
"01101110", 
"01111111", 
"10011110", 
"10000001", 
"01110100", 
"10100010", 
"01011000", 
"01101111", 
"10111101", 
"11001101", 
"01111000", 
"01110010", 
"01111010", 
"10100101", 
"01111011", 
"10110011", 
"01111110", 
"01111001", 
"10001000", 
"01110111", 
"10001000", 
"01010101", 
"01000101", 
"10001010", 
"01100100", 
"10000011", 
"01101100", 
"10001011", 
"10001101", 
"01111110", 
"01101000", 
"01011001", 
"01111100", 
"10110000", 
"10010011", 
"01010110", 
"10001110", 
"01100111", 
"10010110", 
"01000110", 
"01001111", 
"01111110", 
"01110001", 
"10000110", 
"10100101", 
"10101011", 
"01000111", 
"01100011", 
"01101101", 
"10001000", 
"10001101", 
"10010010", 
"01100001", 
"10010100", 
"10100111", 
"10010011", 
"01100011", 
"10010010", 
"10000001", 
"01110100", 
"10001101", 
"01111101", 
"10010100", 
"01011101", 
"10000010", 
"10011010", 
"10011110", 
"10010010", 
"01101011", 
"01100111", 
"10000111", 
"10111110", 
"10011010", 
"01010100", 
"10001000", 
"01111111", 
"10001011", 
"10101000", 
"01110010", 
"10100001", 
"10000011", 
"10101011", 
"10001100", 
"01100111", 
"10001010", 
"10000010", 
"10001011", 
"10001010", 
"10101011", 
"01101110", 
"10001001", 
"01111110", 
"10011000", 
"10011101", 
"10000001", 
"01101000", 
"01111001", 
"10110000", 
"10011001", 
"10110101", 
"01101100", 
"01100101", 
"01111101", 
"01011101", 
"10000010", 
"10000111", 
"10001010", 
"10001001", 
"10000001", 
"01110001", 
"01011010", 
"01101110", 
"10001100", 
"10101101", 
"10010100", 
"10011101", 
"01100100", 
"01100110", 
"10100001", 
"10000000", 
"01100001", 
"11000110", 
"01111001", 
"01101010", 
"10010110", 
"01101100", 
"01101101", 
"01111101", 
"01110101", 
"10010001", 
"10111111", 
"01110101", 
"10010000", 
"01100001", 
"01110110", 
"01010010", 
"10000001", 
"01101001", 
"01111011", 
"10001000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_21: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_21(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
