use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_74_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_74_LAYER;

architecture Behavioral of ROM_FC_84_74_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_74: ROM_ARRAY_PESOS_FC_84 := (
"01011000", 
"01010110", 
"01110100", 
"01101011", 
"10011010", 
"10010010", 
"01111000", 
"01011011", 
"01101101", 
"10101010", 
"01110001", 
"10001100", 
"10010001", 
"01101101", 
"01010100", 
"10010000", 
"10000101", 
"10001111", 
"01110100", 
"10001000", 
"01011110", 
"01100011", 
"01110001", 
"01101000", 
"01101111", 
"10010000", 
"10000001", 
"10011010", 
"01110100", 
"01011001", 
"10001101", 
"01111000", 
"01100010", 
"10100111", 
"01101011", 
"10001011", 
"01100101", 
"10001010", 
"01101010", 
"01011000", 
"10100010", 
"10100111", 
"10001111", 
"01100111", 
"10001100", 
"01001111", 
"10011001", 
"01111011", 
"01011100", 
"01111110", 
"01011001", 
"10110011", 
"01110011", 
"01111010", 
"01101110", 
"10011111", 
"10001101", 
"10001111", 
"01110010", 
"10001010", 
"01101100", 
"00101001", 
"01100000", 
"01011100", 
"01111010", 
"01111001", 
"10001111", 
"01101110", 
"01101011", 
"01100001", 
"01100111", 
"01010001", 
"01011000", 
"10011000", 
"01101111", 
"10011101", 
"01111110", 
"10000011", 
"10011001", 
"01101111", 
"01111011", 
"10011110", 
"10100010", 
"01101000", 
"10001011", 
"10000010", 
"01111000", 
"01100110", 
"10010100", 
"10001000", 
"10001010", 
"10010001", 
"10010101", 
"01001000", 
"10000110", 
"01111111", 
"10000001", 
"01111110", 
"10011000", 
"01111011", 
"10001010", 
"01011111", 
"10101001", 
"01010111", 
"01100001", 
"01110001", 
"01101010", 
"01110110", 
"10101111", 
"10010101", 
"10011101", 
"10001010", 
"10011100", 
"01111001", 
"10000001", 
"10110010", 
"10001001", 
"01111101", 
"01101101", 
"10001001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_74: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_74(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
