use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_71_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_71_LAYER;

architecture Behavioral of ROM_FC_84_71_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_71: ROM_ARRAY_PESOS_FC_84 := (
"01001100", 
"01101010", 
"10001001", 
"01101110", 
"01111110", 
"10010100", 
"01110110", 
"00111111", 
"01100001", 
"10100000", 
"10010101", 
"10100001", 
"01111010", 
"10010010", 
"01100101", 
"10000111", 
"01110010", 
"01011100", 
"10000011", 
"01100001", 
"10010001", 
"01110011", 
"10001001", 
"10011110", 
"01101101", 
"10011010", 
"01100101", 
"10001000", 
"10000011", 
"10011100", 
"10010010", 
"01111101", 
"10001110", 
"01100100", 
"01110110", 
"01101100", 
"01110011", 
"01011010", 
"01010000", 
"01111011", 
"01110010", 
"01101100", 
"01011110", 
"10001100", 
"01011010", 
"01001101", 
"01101010", 
"10000110", 
"10100010", 
"01111001", 
"10011000", 
"01101001", 
"10000001", 
"10010100", 
"01010111", 
"01110110", 
"10011111", 
"01101110", 
"01110110", 
"01010011", 
"01110111", 
"01111001", 
"10011000", 
"01100010", 
"01101101", 
"01100010", 
"01101001", 
"10000000", 
"01101001", 
"10000111", 
"01101000", 
"01101010", 
"01100001", 
"01000001", 
"10000100", 
"10000001", 
"01011010", 
"10000001", 
"10000001", 
"01111011", 
"01100101", 
"01011111", 
"01000001", 
"01110111", 
"01001011", 
"01101110", 
"01110110", 
"10000101", 
"10000000", 
"01111001", 
"01000110", 
"01110010", 
"01111111", 
"01100010", 
"01000011", 
"01101010", 
"00111001", 
"01100100", 
"01010111", 
"10000100", 
"01101100", 
"01010110", 
"10010101", 
"01111101", 
"01101001", 
"01110011", 
"01101000", 
"01110110", 
"01101101", 
"10011001", 
"01110001", 
"10010101", 
"01111001", 
"01110111", 
"01101100", 
"01110001", 
"10110001", 
"01110001", 
"01110100", 
"01101100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_71: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_71(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
