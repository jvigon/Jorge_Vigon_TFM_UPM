use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_69_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_69_LAYER;

architecture Behavioral of ROM_FC_120_69_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_69: ROM_ARRAY_PESOS_FC_120 := (
"01101111", 
"01101110", 
"10100001", 
"01111011", 
"01111010", 
"01101001", 
"01100111", 
"01000101", 
"10000110", 
"10101000", 
"01100100", 
"10110010", 
"10000010", 
"10001011", 
"01101101", 
"10010111", 
"10000100", 
"10011100", 
"10001100", 
"10011110", 
"01101100", 
"10000101", 
"10001111", 
"01101000", 
"01101101", 
"10010001", 
"10000101", 
"10101001", 
"01110111", 
"01100011", 
"01110100", 
"01111001", 
"01111011", 
"01110001", 
"01111010", 
"01011101", 
"10000010", 
"10101111", 
"01110101", 
"10000001", 
"10001101", 
"10010111", 
"01110101", 
"10001110", 
"10000101", 
"01110110", 
"10011100", 
"01101011", 
"10001011", 
"10000101", 
"01110100", 
"01101001", 
"01111101", 
"10010001", 
"01110101", 
"01011001", 
"10000011", 
"10011111", 
"01100000", 
"01100011", 
"10111100", 
"01001111", 
"01110110", 
"10000100", 
"01101111", 
"10001101", 
"01010100", 
"00110001", 
"01101100", 
"01101100", 
"01110011", 
"10010101", 
"01101100", 
"10101001", 
"01110111", 
"10011110", 
"10000011", 
"01110100", 
"10001110", 
"01110001", 
"01101100", 
"10001101", 
"01001110", 
"01011100", 
"01100111", 
"10010000", 
"01101101", 
"01100000", 
"10010100", 
"10001111", 
"10001001", 
"10010101", 
"10011010", 
"10010011", 
"01111111", 
"01110111", 
"01111100", 
"01111101", 
"01001010", 
"01001001", 
"10000101", 
"10001011", 
"01101101", 
"01110000", 
"01100010", 
"10010110", 
"10001001", 
"01111110", 
"01010111", 
"01111010", 
"01110110", 
"10000001", 
"01110110", 
"01011001", 
"10011000", 
"10011110", 
"10001011", 
"01100011", 
"01101001", 
"01110100", 
"01111101", 
"10010000", 
"10000110", 
"01010010", 
"01001100", 
"01101000", 
"01111011", 
"10001001", 
"01100101", 
"10000100", 
"01110001", 
"00110001", 
"10001111", 
"01101010", 
"01110011", 
"01010101", 
"01100111", 
"01011101", 
"01101000", 
"01110000", 
"10001010", 
"10000011", 
"01110101", 
"10001111", 
"10000011", 
"01110010", 
"10001100", 
"10010101", 
"01110110", 
"10111111", 
"00111101", 
"10001101", 
"10010000", 
"01101101", 
"01111011", 
"01011010", 
"10110101", 
"10001001", 
"01111011", 
"01110011", 
"01010001", 
"01001001", 
"10010101", 
"01110101", 
"10000100", 
"10001000", 
"01001111", 
"01000000", 
"01111110", 
"10001011", 
"10100100", 
"01101100", 
"10001111", 
"01100111", 
"01111101", 
"01100010", 
"01100110", 
"00110011", 
"10101000", 
"01110011", 
"01111111", 
"00110101", 
"01111110", 
"00111100", 
"01101011", 
"10100101", 
"01101100", 
"10100010", 
"10001110", 
"01000001", 
"01101111", 
"01110110", 
"10000011", 
"10100010", 
"01000001", 
"01000000", 
"01101111", 
"10101110", 
"10100101", 
"01001010", 
"01110010", 
"01011110", 
"01100001", 
"11000011", 
"00101000", 
"10001010", 
"10000001", 
"01110100", 
"10000110", 
"10101101", 
"01000100", 
"00111100", 
"01101110", 
"10100110", 
"10011100", 
"01101001", 
"01101001", 
"01010101", 
"10100000", 
"01111110", 
"00111010", 
"01111101", 
"01101101", 
"01110001", 
"01001010", 
"01001110", 
"01000110", 
"01111100", 
"10000010", 
"01100001", 
"10010100", 
"01101100", 
"10000001", 
"10101000", 
"11010001", 
"00110100", 
"10000001", 
"10010011", 
"10001011", 
"01101111", 
"01001111", 
"01110100", 
"01101101", 
"01001011", 
"01110010", 
"01011001", 
"10100100", 
"01101110", 
"01101100", 
"10011000", 
"01110011", 
"10010001", 
"00110010", 
"10010110", 
"01111111", 
"01110000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_69: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_69(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
