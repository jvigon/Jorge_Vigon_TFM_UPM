use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_10_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_10_LAYER;

architecture Behavioral of ROM_FC_120_10_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_10: ROM_ARRAY_PESOS_FC_120 := (
"10001001", 
"01111111", 
"01101101", 
"10001001", 
"01110011", 
"10010110", 
"01010110", 
"10001001", 
"01110010", 
"01100011", 
"01110110", 
"01111010", 
"01000011", 
"01110101", 
"10000011", 
"10001101", 
"01110000", 
"01011110", 
"01111000", 
"10001000", 
"01101100", 
"10000100", 
"01011010", 
"01110101", 
"01100100", 
"01111101", 
"10000010", 
"10000111", 
"01010001", 
"10110000", 
"10001011", 
"01111011", 
"01101111", 
"01010001", 
"01011001", 
"01110001", 
"10001101", 
"01101100", 
"10010010", 
"01111000", 
"01011001", 
"10001110", 
"01110111", 
"01101110", 
"01111100", 
"10110011", 
"01110110", 
"10010001", 
"01111100", 
"01010110", 
"01011000", 
"01101110", 
"01101110", 
"10001100", 
"01101100", 
"01111100", 
"01100010", 
"01111110", 
"01100100", 
"01111000", 
"01110001", 
"10101000", 
"10001111", 
"01110111", 
"01110111", 
"01011001", 
"01100111", 
"10000010", 
"01101101", 
"01111000", 
"01111010", 
"10001000", 
"10001101", 
"01101111", 
"01110001", 
"01110110", 
"10000000", 
"01101010", 
"01101111", 
"10011011", 
"10000010", 
"01010101", 
"10000000", 
"10000110", 
"01110100", 
"01111010", 
"01101101", 
"01111011", 
"01011101", 
"01011111", 
"01111000", 
"01101101", 
"01110101", 
"10100100", 
"10001000", 
"01110100", 
"01010111", 
"01010100", 
"01011000", 
"01101011", 
"01110011", 
"10000100", 
"10100000", 
"01101101", 
"01100000", 
"01100010", 
"01110100", 
"01110011", 
"10010010", 
"10010010", 
"10001010", 
"01110111", 
"01110101", 
"01101000", 
"01111010", 
"01100001", 
"01110000", 
"01110011", 
"01110000", 
"01101101", 
"01101101", 
"01111111", 
"01110011", 
"01111001", 
"01111001", 
"10000111", 
"01110000", 
"10010011", 
"01100100", 
"01100001", 
"01101101", 
"10000010", 
"01110011", 
"01111010", 
"01101110", 
"01100001", 
"10000010", 
"10000111", 
"01111101", 
"01110100", 
"01101101", 
"01100100", 
"10000110", 
"10001110", 
"01011100", 
"10010010", 
"01110011", 
"01111111", 
"01111101", 
"01100100", 
"01111111", 
"01101110", 
"01001111", 
"01110011", 
"01011110", 
"01100100", 
"01010001", 
"10001000", 
"01101100", 
"10011101", 
"01110000", 
"10000101", 
"01011000", 
"10010011", 
"01111011", 
"01101011", 
"10100000", 
"01001110", 
"01111100", 
"01111101", 
"01111101", 
"01011110", 
"01101111", 
"01110101", 
"10001110", 
"10010100", 
"10000001", 
"01110001", 
"01101100", 
"10000001", 
"01101111", 
"01111111", 
"01101101", 
"01101011", 
"01011110", 
"01110001", 
"01100111", 
"01101001", 
"01111110", 
"01110101", 
"10001111", 
"01111111", 
"01110100", 
"01111110", 
"01100110", 
"10001101", 
"10001101", 
"01100001", 
"01101011", 
"01110100", 
"01110001", 
"01011110", 
"10011000", 
"01110011", 
"01011011", 
"01111100", 
"10000111", 
"01111100", 
"01100000", 
"10001011", 
"01101000", 
"01100000", 
"10001010", 
"01111000", 
"01111100", 
"01101110", 
"10000000", 
"01110010", 
"01100111", 
"01001101", 
"01101100", 
"10001110", 
"01110011", 
"10000100", 
"01111101", 
"01111010", 
"01100100", 
"10000100", 
"10000000", 
"10001100", 
"01111110", 
"10000100", 
"10000001", 
"01101101", 
"01111100", 
"01010111", 
"10000011", 
"01111100", 
"10010001", 
"01110111", 
"01110010", 
"01111001", 
"01111000", 
"10001111", 
"10000100", 
"01110111", 
"01111101", 
"01110001", 
"01110011", 
"01110011", 
"01101101", 
"01110111", 
"01100100", 
"10010000", 
"10001101", 
"01111011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_10: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_10(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
