use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_72_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_72_LAYER;

architecture Behavioral of ROM_FC_84_72_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_72: ROM_ARRAY_PESOS_FC_84 := (
"10101010", 
"10000010", 
"01100100", 
"10000001", 
"10000010", 
"01111101", 
"01101011", 
"01010101", 
"10000011", 
"01100100", 
"01110000", 
"01111010", 
"01101101", 
"01110010", 
"01101111", 
"01110001", 
"01110110", 
"01100111", 
"01111001", 
"01101111", 
"01111110", 
"01001101", 
"01010111", 
"01101110", 
"01100010", 
"10010001", 
"01000110", 
"01110001", 
"01010110", 
"01100111", 
"01110001", 
"10101010", 
"10000001", 
"01010010", 
"01011010", 
"00100000", 
"10011001", 
"01111010", 
"10110010", 
"01100110", 
"10010011", 
"11000010", 
"10010100", 
"01001101", 
"01010100", 
"01110000", 
"01010000", 
"10000000", 
"10000110", 
"01110110", 
"01001010", 
"10001010", 
"01101101", 
"01101011", 
"10000111", 
"10000110", 
"10011011", 
"10000001", 
"01011111", 
"01010010", 
"01111010", 
"10000000", 
"01010001", 
"01100101", 
"01100010", 
"00111111", 
"10001000", 
"01110100", 
"01100110", 
"01110000", 
"10001100", 
"10001011", 
"01001100", 
"01111100", 
"10100101", 
"10010111", 
"10000011", 
"01111110", 
"10000101", 
"01110001", 
"01110011", 
"10011000", 
"01111100", 
"10011100", 
"01110111", 
"01101101", 
"01100001", 
"10000100", 
"01110001", 
"10100101", 
"10010001", 
"01101101", 
"10010011", 
"01001001", 
"01101111", 
"10100100", 
"10000011", 
"01111111", 
"10001110", 
"10001001", 
"10000011", 
"10001100", 
"10010101", 
"01001001", 
"01000001", 
"10000011", 
"01101000", 
"01110110", 
"10000110", 
"01111000", 
"01011000", 
"10001100", 
"01101101", 
"01101110", 
"01100000", 
"01110111", 
"10010111", 
"00011001", 
"10010001", 
"01100010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_72: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_72(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
