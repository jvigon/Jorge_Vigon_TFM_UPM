use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_21_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_21_LAYER;

architecture Behavioral of ROM_FC_84_21_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_21: ROM_ARRAY_PESOS_FC_84 := (
"01111000", 
"01100000", 
"01100001", 
"10001000", 
"10100100", 
"10001110", 
"10001000", 
"01011011", 
"01110101", 
"10100101", 
"01110100", 
"10001101", 
"01001101", 
"01100110", 
"01001011", 
"01111000", 
"01100110", 
"10011100", 
"10100000", 
"01110111", 
"10001100", 
"10000010", 
"01111000", 
"01000011", 
"01100111", 
"01000100", 
"10001111", 
"10001101", 
"10100111", 
"01110101", 
"10000101", 
"01111110", 
"10011100", 
"10000010", 
"01101101", 
"01111111", 
"10000001", 
"01111101", 
"01110011", 
"01011110", 
"10000100", 
"01110000", 
"10100010", 
"01100110", 
"01110011", 
"01110101", 
"01101100", 
"01110110", 
"01110101", 
"01100101", 
"01111000", 
"10011000", 
"10000110", 
"01101001", 
"01101101", 
"10100101", 
"10010000", 
"10010100", 
"01111011", 
"01100101", 
"01100111", 
"01110011", 
"01110010", 
"10011100", 
"01101110", 
"01011101", 
"01111000", 
"10000001", 
"01101111", 
"01011110", 
"01111011", 
"10000001", 
"01111000", 
"10100111", 
"10010000", 
"10010010", 
"10011110", 
"10001101", 
"10001000", 
"01110000", 
"10010010", 
"10001000", 
"01111001", 
"01100010", 
"10010010", 
"10001110", 
"01110111", 
"10001100", 
"01101001", 
"01101001", 
"01010101", 
"11000110", 
"01011101", 
"01111111", 
"01011100", 
"01101010", 
"01111011", 
"10000000", 
"01101101", 
"01011111", 
"01100010", 
"01101000", 
"01110000", 
"01100110", 
"10001111", 
"10001101", 
"10001110", 
"01111110", 
"01111111", 
"01100110", 
"10101001", 
"10000010", 
"01111000", 
"01111111", 
"10000100", 
"01110010", 
"01011011", 
"10000100", 
"01100001", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_21 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_21(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
