use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_76_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_76_LAYER;

architecture Behavioral of ROM_FC_120_76_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_76: ROM_ARRAY_PESOS_FC_120 := (
"01101010", 
"10000010", 
"10000110", 
"10100010", 
"10011101", 
"01011110", 
"01110110", 
"01110101", 
"10001110", 
"10100101", 
"10110100", 
"10010000", 
"10010101", 
"11110100", 
"10001101", 
"01101011", 
"01011000", 
"01110000", 
"10101010", 
"10011010", 
"01111110", 
"01110101", 
"01010010", 
"01110111", 
"10001101", 
"10001010", 
"01110110", 
"10001010", 
"10000010", 
"10001100", 
"01101011", 
"10001100", 
"01100111", 
"10011101", 
"01011001", 
"01111010", 
"10001010", 
"01110101", 
"01101110", 
"01111001", 
"10000010", 
"01110001", 
"01101100", 
"10001100", 
"01110000", 
"10110111", 
"01110001", 
"01111011", 
"01111110", 
"01111101", 
"10101011", 
"01100110", 
"01111111", 
"01100101", 
"01100010", 
"10001110", 
"01101011", 
"01011011", 
"01011100", 
"01110110", 
"01110111", 
"10000110", 
"01110001", 
"01111101", 
"01111000", 
"01101100", 
"01110111", 
"01000000", 
"01101111", 
"01111010", 
"01000110", 
"01100100", 
"01110000", 
"01101010", 
"10010111", 
"10001011", 
"10011000", 
"01100101", 
"10001100", 
"01101010", 
"01101101", 
"10101011", 
"10001011", 
"01101011", 
"10000110", 
"10000001", 
"10000001", 
"01111000", 
"01101011", 
"10010111", 
"10001011", 
"01110111", 
"01110001", 
"00111001", 
"01111010", 
"10001100", 
"10001011", 
"10001111", 
"01100101", 
"01110100", 
"01111101", 
"01011011", 
"01101111", 
"10101001", 
"01101111", 
"01101111", 
"01100101", 
"01101010", 
"01111000", 
"00001000", 
"10001110", 
"01110010", 
"10000111", 
"10001000", 
"10001011", 
"01100101", 
"01111110", 
"00111100", 
"01011001", 
"01111100", 
"01110010", 
"10010001", 
"10001100", 
"01011110", 
"01111011", 
"01011101", 
"10000000", 
"10000000", 
"01101011", 
"01011011", 
"01101100", 
"01001100", 
"01100010", 
"01010110", 
"00001001", 
"01011111", 
"01110100", 
"10011000", 
"01111111", 
"10001010", 
"01100010", 
"01100001", 
"01101010", 
"01101000", 
"01000001", 
"00111010", 
"01010110", 
"01011101", 
"10000001", 
"01111001", 
"00110100", 
"01101000", 
"01011001", 
"10011011", 
"10010001", 
"10010100", 
"10010000", 
"00110011", 
"10001110", 
"10001111", 
"10000100", 
"01100010", 
"10010110", 
"10100001", 
"10000101", 
"01111000", 
"00111101", 
"10100101", 
"01110010", 
"10001010", 
"01100101", 
"01110000", 
"01111101", 
"11001111", 
"01101110", 
"10001001", 
"10000000", 
"10001100", 
"01101101", 
"01110100", 
"10000111", 
"01011111", 
"01110100", 
"10100111", 
"01101111", 
"01000000", 
"00101111", 
"01100011", 
"10000000", 
"01110100", 
"10000010", 
"01110111", 
"10001001", 
"10011001", 
"00110100", 
"00011101", 
"01111001", 
"01110010", 
"01101100", 
"01101001", 
"10001001", 
"01010111", 
"01100001", 
"10010010", 
"10010010", 
"10110100", 
"01111001", 
"10001010", 
"00111101", 
"10011010", 
"01110100", 
"00101110", 
"01101001", 
"01011001", 
"10011110", 
"01000010", 
"10000000", 
"10001010", 
"00101100", 
"01110011", 
"11000010", 
"10011010", 
"01111110", 
"10000000", 
"01101110", 
"11000011", 
"01110010", 
"01101001", 
"01111000", 
"01110010", 
"01100000", 
"10000010", 
"10001100", 
"01001100", 
"01011100", 
"01111011", 
"11011011", 
"10101101", 
"01111011", 
"10001000", 
"10010000", 
"10110110", 
"00111100", 
"01110110", 
"10001101", 
"10001111", 
"10000111", 
"01110011", 
"10001010", 
"01001101", 
"01000100", 
"01011100", 
"10100111", 
"10111011", 
"01101100", 
"01100111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_76: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_76(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
