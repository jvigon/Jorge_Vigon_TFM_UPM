use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_14_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_14_LAYER;

architecture Behavioral of ROM_FC_120_14_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_14: ROM_ARRAY_PESOS_FC_120 := (
"11000000", 
"10110000", 
"10011000", 
"10011001", 
"01011000", 
"10101000", 
"01100111", 
"10000101", 
"10110100", 
"01110011", 
"11010110", 
"01111100", 
"01111000", 
"11111000", 
"10101000", 
"01100010", 
"10101001", 
"10110100", 
"01010010", 
"00110001", 
"01110001", 
"01111101", 
"10010110", 
"01100011", 
"01011101", 
"10001011", 
"01111110", 
"00110111", 
"01111011", 
"10101100", 
"10001000", 
"01000110", 
"01001011", 
"01110011", 
"00010100", 
"00101011", 
"01111101", 
"01111101", 
"10000000", 
"01001011", 
"01110010", 
"01100110", 
"01111010", 
"01110110", 
"01011100", 
"00100010", 
"10000000", 
"01010011", 
"01100011", 
"00000000", 
"01111000", 
"10100001", 
"10011001", 
"10101000", 
"10101100", 
"01110001", 
"10111101", 
"01110000", 
"10001010", 
"01011110", 
"01011010", 
"01101110", 
"10001110", 
"01110100", 
"01101000", 
"00110010", 
"01101100", 
"10111011", 
"01011100", 
"01100010", 
"10101100", 
"01101100", 
"10101100", 
"10000100", 
"11010011", 
"01011010", 
"10011101", 
"10101000", 
"01111001", 
"10001001", 
"10010101", 
"01101011", 
"01110001", 
"01101110", 
"10110010", 
"01110001", 
"01101111", 
"10100100", 
"10101001", 
"10000011", 
"01100111", 
"01011100", 
"01111011", 
"10101010", 
"01110001", 
"01110011", 
"01111110", 
"01101011", 
"10010101", 
"01101110", 
"01101110", 
"01110000", 
"01111001", 
"01101010", 
"10011011", 
"01011000", 
"01011111", 
"01111011", 
"10010101", 
"10001100", 
"01111010", 
"01110110", 
"01000010", 
"01000100", 
"00011101", 
"01000101", 
"10000101", 
"10001000", 
"10000111", 
"00100110", 
"11000010", 
"01101101", 
"10000001", 
"01100000", 
"01111110", 
"01001000", 
"01111101", 
"10100110", 
"10101011", 
"10100100", 
"00111011", 
"01010100", 
"01101001", 
"10010001", 
"01110110", 
"10000011", 
"01101010", 
"11000011", 
"11011000", 
"01110010", 
"01100001", 
"10000111", 
"01111011", 
"01110001", 
"01110100", 
"10001110", 
"01100100", 
"01100110", 
"01111111", 
"10101001", 
"01101011", 
"01110111", 
"01101010", 
"10001000", 
"10011010", 
"01010100", 
"10010100", 
"01100100", 
"10001001", 
"10100010", 
"01110011", 
"10001110", 
"01100110", 
"00111011", 
"01110001", 
"01000010", 
"01011000", 
"01101100", 
"01110100", 
"10001000", 
"01001100", 
"01111011", 
"10100111", 
"10011010", 
"01110101", 
"10001011", 
"01011100", 
"10110011", 
"01100000", 
"00101011", 
"01111111", 
"10000001", 
"01111010", 
"00010110", 
"10011000", 
"01000010", 
"01001110", 
"01111001", 
"10001010", 
"01110010", 
"10001100", 
"10011011", 
"01110011", 
"01001111", 
"01000011", 
"01010010", 
"01101101", 
"01111011", 
"01101000", 
"01110110", 
"01100110", 
"10001110", 
"01101110", 
"10001010", 
"01010111", 
"01110100", 
"10000010", 
"01111100", 
"10001111", 
"10011100", 
"01111011", 
"10000000", 
"10000000", 
"10011010", 
"00110000", 
"01010011", 
"10001001", 
"10000000", 
"10011000", 
"10000111", 
"01100000", 
"01010111", 
"01100101", 
"01111010", 
"01111101", 
"10010010", 
"01100011", 
"01111000", 
"01011101", 
"01101100", 
"01011111", 
"00011010", 
"10001111", 
"01011110", 
"10001100", 
"10101101", 
"01011100", 
"10100011", 
"01101111", 
"10001101", 
"01101111", 
"01110001", 
"00110000", 
"01000100", 
"01110100", 
"01000011", 
"10000011", 
"01011001", 
"01111100", 
"01111111", 
"01100101", 
"01110011", 
"01110100", 
"10000101", 
"10000010", 
"10001100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_14: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_14(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
