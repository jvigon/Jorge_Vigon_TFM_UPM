use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_79_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_79_LAYER;

architecture Behavioral of ROM_FC_120_79_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_79: ROM_ARRAY_PESOS_FC_120 := (
"01101010", 
"01111111", 
"10011110", 
"01101110", 
"10010001", 
"00110101", 
"10011111", 
"10001000", 
"10001000", 
"01010110", 
"01011110", 
"01010110", 
"10100110", 
"01110110", 
"10000110", 
"01011011", 
"01111000", 
"01101001", 
"10000110", 
"00101111", 
"01111010", 
"01011101", 
"01110100", 
"01100100", 
"10001111", 
"01101001", 
"01100100", 
"01110010", 
"10000010", 
"10000000", 
"10000010", 
"01111111", 
"01101100", 
"01010101", 
"10001010", 
"01101100", 
"10001000", 
"01111111", 
"01101101", 
"01011101", 
"01110100", 
"10000010", 
"10000111", 
"01110010", 
"10000100", 
"10100000", 
"01111111", 
"01110011", 
"01101100", 
"01101111", 
"01101101", 
"10001111", 
"01111000", 
"01110011", 
"01111100", 
"01001010", 
"01111010", 
"01011010", 
"01111001", 
"10001010", 
"01110000", 
"01110010", 
"01110000", 
"01110011", 
"01111011", 
"10001100", 
"10010010", 
"10010110", 
"01111101", 
"10101100", 
"01100101", 
"01111001", 
"01110011", 
"01110110", 
"10101010", 
"01011011", 
"01110001", 
"01000010", 
"10000111", 
"10001000", 
"10001011", 
"10000101", 
"10001000", 
"01001110", 
"10001010", 
"01100111", 
"01011111", 
"01101100", 
"01111000", 
"01110010", 
"10010010", 
"01011110", 
"01000011", 
"01100000", 
"01110100", 
"01111000", 
"01111101", 
"01111000", 
"10000010", 
"01001000", 
"01111000", 
"01110111", 
"01100101", 
"01100100", 
"01110110", 
"10001000", 
"01010000", 
"10001111", 
"00010100", 
"01110100", 
"01111000", 
"01100100", 
"01100011", 
"10001000", 
"01001111", 
"01100011", 
"01111011", 
"10000011", 
"10110100", 
"01100101", 
"10000101", 
"01100100", 
"01111011", 
"10001101", 
"01000110", 
"01001110", 
"10000111", 
"01110001", 
"10100101", 
"01101010", 
"01100101", 
"10101010", 
"01110110", 
"10110001", 
"01000000", 
"01111110", 
"10000111", 
"01110010", 
"10111011", 
"01100010", 
"00111001", 
"01100000", 
"10000010", 
"01101011", 
"10000000", 
"01110110", 
"10000101", 
"10000100", 
"10001101", 
"01110110", 
"01111010", 
"10101011", 
"10010101", 
"01100001", 
"01110101", 
"01001111", 
"01010100", 
"10001100", 
"01110000", 
"01111101", 
"01011111", 
"01101000", 
"01100001", 
"01001000", 
"10001010", 
"10001110", 
"10001110", 
"10001101", 
"10001000", 
"01001101", 
"01110110", 
"10010000", 
"10000111", 
"10011110", 
"10000010", 
"10011001", 
"01111101", 
"01111010", 
"01101011", 
"01011100", 
"01110000", 
"01101010", 
"10011000", 
"01111000", 
"01110101", 
"01010110", 
"01100101", 
"01111011", 
"10000111", 
"01110110", 
"01110111", 
"10010110", 
"10000011", 
"01101100", 
"10001011", 
"10010110", 
"10001011", 
"10101000", 
"01100111", 
"01111011", 
"10000101", 
"01101001", 
"10101011", 
"01101011", 
"01010001", 
"10010010", 
"10000000", 
"01111000", 
"10000011", 
"10000000", 
"10001101", 
"10011101", 
"10000100", 
"01011001", 
"10011000", 
"01110111", 
"01110011", 
"01111001", 
"01011100", 
"01101101", 
"01011000", 
"10010010", 
"10000110", 
"01110010", 
"01111011", 
"01011111", 
"01101001", 
"01111010", 
"01111001", 
"01101011", 
"10101011", 
"01101100", 
"10001110", 
"01110111", 
"01010111", 
"01110110", 
"10100100", 
"01110010", 
"10000000", 
"01110100", 
"10010011", 
"01100111", 
"01110000", 
"01010011", 
"10001011", 
"01111100", 
"10011101", 
"10001000", 
"10000110", 
"10010001", 
"01010101", 
"01011111", 
"11000000", 
"01100000", 
"10010101", 
"10001111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_79: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_79(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
