use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_35_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_35_LAYER;

architecture Behavioral of ROM_FC_120_35_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_35: ROM_ARRAY_PESOS_FC_120 := (
"01011111", 
"01000001", 
"01100011", 
"10110110", 
"10011011", 
"10000011", 
"10010011", 
"01011111", 
"10001001", 
"10011100", 
"10100011", 
"00100000", 
"10011100", 
"01100011", 
"10001010", 
"10000001", 
"01111000", 
"10000111", 
"10101001", 
"10110100", 
"10010110", 
"00011111", 
"10010011", 
"01111011", 
"01110011", 
"01101011", 
"01111010", 
"01111100", 
"01110001", 
"01111100", 
"10000111", 
"01100101", 
"01110010", 
"10101111", 
"10100101", 
"10011010", 
"10001110", 
"01110000", 
"01010001", 
"01101010", 
"10000101", 
"01111101", 
"01111111", 
"01110001", 
"10000110", 
"10100111", 
"01111011", 
"01011110", 
"10010110", 
"10101110", 
"01111101", 
"01101101", 
"01111111", 
"01001111", 
"01000111", 
"01110100", 
"01110110", 
"01111011", 
"01111101", 
"10010011", 
"01010101", 
"10100101", 
"01111000", 
"10000011", 
"10000011", 
"10011001", 
"10101011", 
"11101100", 
"10001100", 
"01011010", 
"10011111", 
"01011010", 
"01111011", 
"00110111", 
"10011010", 
"01001101", 
"01000011", 
"10000000", 
"01110000", 
"01111100", 
"01001101", 
"01111000", 
"10000100", 
"11100100", 
"10000111", 
"00101001", 
"10001101", 
"01010101", 
"10001110", 
"01011010", 
"01111111", 
"01001000", 
"10000110", 
"01110001", 
"01110011", 
"01110111", 
"01111011", 
"10001101", 
"10001101", 
"10011000", 
"01101100", 
"10010001", 
"01110001", 
"01011111", 
"10010001", 
"01101001", 
"01110110", 
"01100001", 
"10010011", 
"01100111", 
"01111010", 
"10001110", 
"10000101", 
"10011010", 
"10001111", 
"01100011", 
"01100101", 
"10010101", 
"01100100", 
"10001110", 
"01110111", 
"10001001", 
"01111101", 
"01100010", 
"10001011", 
"01110110", 
"01111100", 
"01111110", 
"10010000", 
"11001010", 
"00100101", 
"01110111", 
"10000010", 
"01011001", 
"10100100", 
"01000101", 
"01110110", 
"01111011", 
"01111010", 
"10011010", 
"01111111", 
"01101110", 
"01111111", 
"10000011", 
"01001111", 
"10100111", 
"01011010", 
"10010101", 
"01111101", 
"01100000", 
"01111111", 
"01111100", 
"10000011", 
"10000000", 
"10001001", 
"10010100", 
"01111010", 
"10001110", 
"10000110", 
"01110011", 
"01101011", 
"01110110", 
"10000100", 
"01110111", 
"01110110", 
"10100011", 
"01011100", 
"10010001", 
"01110000", 
"01111010", 
"10000011", 
"10001111", 
"01111110", 
"01110111", 
"10010001", 
"01110010", 
"01100101", 
"01010111", 
"01100101", 
"10000011", 
"10000110", 
"01111011", 
"10001111", 
"01110111", 
"01110000", 
"01110010", 
"01111000", 
"01110000", 
"00000010", 
"10100000", 
"01111111", 
"10000010", 
"10001010", 
"10010111", 
"01011010", 
"10100101", 
"10010101", 
"01011000", 
"01110100", 
"01110011", 
"10000110", 
"01000011", 
"01101100", 
"10010011", 
"01110010", 
"01010111", 
"10000000", 
"10000000", 
"01011100", 
"10011001", 
"10001011", 
"10010110", 
"10000010", 
"01111111", 
"01001111", 
"01011001", 
"10010001", 
"01010011", 
"10001000", 
"01010111", 
"01011010", 
"10010100", 
"10000110", 
"10010011", 
"01100110", 
"01110010", 
"10101110", 
"10010110", 
"01101111", 
"01111111", 
"10001001", 
"01101011", 
"01111101", 
"01100010", 
"01110111", 
"01111011", 
"01100001", 
"01110111", 
"01101100", 
"01111010", 
"10100011", 
"10100011", 
"10100010", 
"10010110", 
"01110110", 
"10011101", 
"10011010", 
"01110101", 
"10000111", 
"01011000", 
"01111100", 
"10011011", 
"10101000", 
"10100100", 
"10000111", 
"10011001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_35: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_35(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
