use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_49_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_49_LAYER;

architecture Behavioral of ROM_FC_84_49_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_49: ROM_ARRAY_PESOS_FC_84 := (
"01111000", 
"01011000", 
"01100000", 
"10000101", 
"10011011", 
"01110101", 
"10000111", 
"10000000", 
"01100101", 
"10100001", 
"10000011", 
"01110011", 
"01011111", 
"10001011", 
"10011000", 
"01100101", 
"01101000", 
"10000000", 
"10000010", 
"01111101", 
"10010011", 
"10100101", 
"10000110", 
"01011100", 
"10010010", 
"10001011", 
"01100001", 
"01100100", 
"01100101", 
"10000101", 
"10001011", 
"10000111", 
"01110101", 
"10010111", 
"01010100", 
"01001110", 
"01111010", 
"01011101", 
"10101111", 
"01100000", 
"00100111", 
"10101100", 
"10001011", 
"10001101", 
"10000011", 
"01010100", 
"01111111", 
"10001100", 
"10101110", 
"01101011", 
"10000101", 
"10110001", 
"10001001", 
"01010100", 
"10001000", 
"10000001", 
"01101111", 
"01101001", 
"01100011", 
"10011110", 
"10011011", 
"10011111", 
"10011001", 
"11000001", 
"01111000", 
"00111011", 
"10010000", 
"10001011", 
"01111110", 
"01110000", 
"01100010", 
"01111111", 
"01010000", 
"01110111", 
"01110001", 
"10000001", 
"10000001", 
"10000111", 
"10010000", 
"01100101", 
"01101100", 
"01101001", 
"01101000", 
"01111111", 
"01111001", 
"10000001", 
"10001111", 
"10001000", 
"10010011", 
"01010100", 
"01111111", 
"10001110", 
"01101100", 
"01101011", 
"01110000", 
"01100110", 
"01001001", 
"01111001", 
"10001011", 
"01111010", 
"01100111", 
"01110111", 
"01001011", 
"10000000", 
"01101111", 
"10000011", 
"10000000", 
"10001110", 
"01110101", 
"00110111", 
"01101100", 
"01011111", 
"10010010", 
"01110011", 
"10000111", 
"01011101", 
"01001010", 
"10011101", 
"01110101", 
"01010101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_49: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_49(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
