use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_76_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_76_LAYER;

architecture Behavioral of ROM_FC_84_76_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_76: ROM_ARRAY_PESOS_FC_84 := (
"01011100", 
"01110111", 
"01100111", 
"10000010", 
"10100011", 
"10001110", 
"10010101", 
"01101000", 
"10011010", 
"10000111", 
"10011000", 
"01111010", 
"01011110", 
"10000111", 
"10111111", 
"01110011", 
"10001000", 
"10001100", 
"01101111", 
"10010101", 
"01101100", 
"01010110", 
"01100111", 
"10000100", 
"01110011", 
"10001100", 
"01110101", 
"01110100", 
"10010010", 
"01101110", 
"10000101", 
"01001100", 
"01101101", 
"10010111", 
"01110111", 
"01011111", 
"10100011", 
"01011110", 
"01110101", 
"01101111", 
"01011111", 
"01110001", 
"10000000", 
"10000110", 
"01010000", 
"01100010", 
"10000100", 
"10011110", 
"10001011", 
"10011101", 
"01110010", 
"10100000", 
"01101111", 
"01100101", 
"10010011", 
"10001101", 
"01101110", 
"01110100", 
"10001000", 
"10011011", 
"01111001", 
"10000011", 
"10011001", 
"01110010", 
"10000101", 
"10000000", 
"01100100", 
"01100001", 
"10000111", 
"10111100", 
"01010001", 
"01100011", 
"01000010", 
"01011110", 
"01101111", 
"01111011", 
"10010000", 
"01111011", 
"01010111", 
"10000011", 
"01111011", 
"10000100", 
"01111110", 
"01110001", 
"01101001", 
"10000100", 
"10011001", 
"01011000", 
"10000101", 
"01010101", 
"00110100", 
"10000000", 
"01101101", 
"01111010", 
"01101010", 
"10000101", 
"01011000", 
"10001101", 
"10000110", 
"01110100", 
"01101111", 
"01110110", 
"01100100", 
"10000000", 
"00111011", 
"10001110", 
"10010001", 
"10001111", 
"01111100", 
"10011101", 
"01111111", 
"01101101", 
"10010111", 
"01011001", 
"01101001", 
"10000100", 
"01110010", 
"01111101", 
"10011100", 
"01011111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_76: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_76(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
