use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_61_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_61_LAYER;

architecture Behavioral of ROM_FC_120_61_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_61: ROM_ARRAY_PESOS_FC_120 := (
"10000011", 
"01111101", 
"10000000", 
"10000101", 
"10001010", 
"10011101", 
"10000011", 
"10000110", 
"10010000", 
"10001001", 
"01011001", 
"01010101", 
"01100101", 
"10010100", 
"10000011", 
"10001001", 
"10011011", 
"10000010", 
"00111011", 
"10000001", 
"10010010", 
"10100100", 
"10011000", 
"11001101", 
"10000010", 
"10010001", 
"01110100", 
"01011011", 
"01011110", 
"01011111", 
"10100000", 
"01111011", 
"10011001", 
"00111010", 
"01010001", 
"01101001", 
"10000101", 
"10011010", 
"10010100", 
"10111100", 
"10010010", 
"10000000", 
"10000101", 
"01111001", 
"01010000", 
"00001001", 
"10000000", 
"10000001", 
"01010001", 
"00111110", 
"01111000", 
"01100001", 
"01110111", 
"01000011", 
"01111011", 
"10011010", 
"01111100", 
"10100100", 
"01101000", 
"01010101", 
"10000110", 
"00000000", 
"01111101", 
"01100010", 
"10010111", 
"01010110", 
"01100011", 
"10000101", 
"01110110", 
"01100111", 
"01000110", 
"10011100", 
"10100010", 
"10110011", 
"10011101", 
"01110010", 
"01101001", 
"10110000", 
"01100110", 
"01101010", 
"01110110", 
"00101001", 
"01100111", 
"01111111", 
"10100101", 
"10000000", 
"10010001", 
"10011001", 
"01101011", 
"10010001", 
"10001011", 
"10011011", 
"10010111", 
"01111110", 
"01111010", 
"01011101", 
"10010110", 
"01001110", 
"01111101", 
"01010101", 
"10100100", 
"10011100", 
"10000000", 
"10010001", 
"10001011", 
"10100101", 
"01011100", 
"00110100", 
"10010000", 
"10011010", 
"01110111", 
"01110100", 
"01010010", 
"01010111", 
"10110011", 
"01100111", 
"10110101", 
"00110111", 
"10000101", 
"10000001", 
"10000101", 
"01111011", 
"00111001", 
"01100101", 
"10011001", 
"10111111", 
"10100000", 
"10001001", 
"01011100", 
"10000011", 
"10010100", 
"01100001", 
"01100111", 
"10000110", 
"01011010", 
"10101011", 
"10001010", 
"10000011", 
"01110111", 
"01011101", 
"10001011", 
"10001001", 
"01110100", 
"01111011", 
"01110011", 
"01011101", 
"10000001", 
"01101100", 
"10100110", 
"01111001", 
"01011101", 
"01111011", 
"10000010", 
"10000100", 
"10000100", 
"01110000", 
"10000110", 
"10001100", 
"01101101", 
"10001110", 
"10001101", 
"10010100", 
"01110001", 
"10011101", 
"10010011", 
"10110110", 
"01010101", 
"01101101", 
"10110011", 
"10011011", 
"01110010", 
"01101101", 
"10011100", 
"10001110", 
"01101110", 
"10000111", 
"01100001", 
"10010111", 
"11000001", 
"10010011", 
"10001000", 
"01010110", 
"01010110", 
"01101100", 
"10011001", 
"01101000", 
"01111110", 
"01101110", 
"10001100", 
"10001000", 
"10010111", 
"01111100", 
"10011101", 
"10010011", 
"01110100", 
"01100111", 
"01110110", 
"10000000", 
"01011011", 
"01110100", 
"01101000", 
"01110010", 
"01110011", 
"01111111", 
"11000110", 
"01101100", 
"01100000", 
"01110111", 
"10001011", 
"01110001", 
"10011000", 
"01100000", 
"01111010", 
"01110110", 
"01101111", 
"10111110", 
"01110011", 
"10011011", 
"01000011", 
"01111000", 
"10100110", 
"01011000", 
"01110111", 
"01111000", 
"01111010", 
"01101011", 
"10010111", 
"10011111", 
"10010001", 
"01111011", 
"10001010", 
"10001011", 
"01110011", 
"10000100", 
"01111110", 
"01101010", 
"01111010", 
"10011111", 
"10001010", 
"01110001", 
"01011111", 
"10010000", 
"11000101", 
"10101011", 
"01101100", 
"01011111", 
"01011110", 
"01001110", 
"01110100", 
"01111111", 
"10000110", 
"01111110", 
"10000111", 
"01110000", 
"01111001", 
"01110100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_61: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_61(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
