use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_78_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_78_LAYER;

architecture Behavioral of ROM_FC_120_78_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_78: ROM_ARRAY_PESOS_FC_120 := (
"10001010", 
"10011001", 
"01110010", 
"10001000", 
"10001011", 
"10010011", 
"01011001", 
"10000000", 
"10001010", 
"00110111", 
"10000011", 
"01111101", 
"01010110", 
"01110001", 
"01101001", 
"10000001", 
"01111011", 
"01100110", 
"01101000", 
"10000100", 
"01101011", 
"01101010", 
"10000101", 
"01110111", 
"01101111", 
"00111011", 
"10001100", 
"01011100", 
"01101010", 
"01111010", 
"01101100", 
"01011110", 
"01001100", 
"10010010", 
"10010010", 
"10100111", 
"10000110", 
"01100101", 
"10001011", 
"10001110", 
"01101111", 
"10000011", 
"10100001", 
"00100000", 
"10000101", 
"10010001", 
"01110000", 
"10000010", 
"01111111", 
"10011000", 
"01111110", 
"01110001", 
"10010010", 
"10001010", 
"01101111", 
"01110101", 
"10010000", 
"10000100", 
"01111111", 
"01110111", 
"01100111", 
"01110110", 
"01111110", 
"01101111", 
"10000110", 
"10101011", 
"10001110", 
"10100111", 
"01100010", 
"01110000", 
"10001011", 
"01100011", 
"10000011", 
"01000000", 
"01010010", 
"10001110", 
"11000011", 
"01101111", 
"01111000", 
"01111110", 
"01100110", 
"10001010", 
"10011110", 
"01101001", 
"01101010", 
"10000111", 
"01110110", 
"01010001", 
"01101100", 
"01010001", 
"01011001", 
"01101000", 
"10011111", 
"01000100", 
"10000111", 
"10000110", 
"01100001", 
"10010111", 
"01111010", 
"10010001", 
"10000111", 
"10001101", 
"10000111", 
"01111101", 
"01111001", 
"01110011", 
"10011011", 
"01010110", 
"01111100", 
"10001101", 
"01111101", 
"10000101", 
"01101011", 
"01110110", 
"01001100", 
"01011111", 
"10001001", 
"10011111", 
"10001110", 
"10000010", 
"10010001", 
"01111100", 
"10001110", 
"01110111", 
"11001111", 
"01010011", 
"01101001", 
"10010010", 
"10010000", 
"10000110", 
"01100110", 
"01000101", 
"01111100", 
"10000011", 
"10011000", 
"01101001", 
"01101011", 
"01111010", 
"01101001", 
"01110111", 
"10010101", 
"00101100", 
"01110001", 
"01101101", 
"01111011", 
"10000001", 
"01110100", 
"00111000", 
"01101010", 
"01100100", 
"01000101", 
"01100110", 
"10000010", 
"01011010", 
"01011101", 
"01010011", 
"01101111", 
"01000110", 
"10000110", 
"01111111", 
"01111111", 
"01011001", 
"01110010", 
"01010111", 
"01110000", 
"10001010", 
"10011101", 
"10001010", 
"01101110", 
"10001000", 
"01111011", 
"01001101", 
"10010010", 
"10010000", 
"10000101", 
"01110010", 
"01111110", 
"01101110", 
"01100110", 
"01110110", 
"01110000", 
"10010001", 
"01011001", 
"01110101", 
"10001000", 
"01010010", 
"10001011", 
"01100110", 
"01100110", 
"10001111", 
"01110101", 
"10001001", 
"01111011", 
"01100100", 
"01111101", 
"10000111", 
"10001010", 
"01110111", 
"01100100", 
"01100010", 
"01111110", 
"01101100", 
"01100101", 
"10001011", 
"10000100", 
"01100000", 
"10001111", 
"10001100", 
"01011100", 
"01110001", 
"10010101", 
"01111001", 
"01101010", 
"01110101", 
"01011000", 
"01111101", 
"10001000", 
"01011000", 
"01011100", 
"01100010", 
"01011111", 
"01100101", 
"01110011", 
"10000010", 
"01011100", 
"01010000", 
"10010110", 
"01110110", 
"10001101", 
"01100110", 
"01010110", 
"10101101", 
"01111010", 
"01100011", 
"01100010", 
"01010001", 
"01111000", 
"01110010", 
"01111011", 
"10001000", 
"10001000", 
"10000010", 
"10000100", 
"10000000", 
"01110110", 
"10011001", 
"10111111", 
"10001110", 
"01110001", 
"01011010", 
"01101101", 
"01101011", 
"01101111", 
"01101000", 
"10000010", 
"10000001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_78: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_78(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
