use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_107_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_107_LAYER;

architecture Behavioral of ROM_FC_120_107_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_107: ROM_ARRAY_PESOS_FC_120 := (
"01111010", 
"10000000", 
"01100100", 
"01101110", 
"10000100", 
"01110100", 
"01101111", 
"01110001", 
"01101111", 
"01100011", 
"01101101", 
"01111011", 
"01110100", 
"01011100", 
"01111011", 
"01101111", 
"01111100", 
"01111001", 
"01100110", 
"01101111", 
"01111010", 
"01100110", 
"01110110", 
"10001000", 
"01111110", 
"01011111", 
"01100010", 
"01111011", 
"10000001", 
"10000100", 
"01111011", 
"10001100", 
"01110100", 
"01110111", 
"10001111", 
"01110110", 
"01101111", 
"01111111", 
"01110110", 
"01011011", 
"10000110", 
"01111001", 
"01111011", 
"10010101", 
"01110100", 
"01101110", 
"10001000", 
"10000101", 
"01110100", 
"01110001", 
"10011110", 
"01100001", 
"10000100", 
"01111111", 
"01100110", 
"10000010", 
"01110010", 
"01111011", 
"10001010", 
"01100000", 
"01100111", 
"01101000", 
"10001111", 
"01111100", 
"01111011", 
"01111001", 
"10000100", 
"10001000", 
"01100101", 
"01111110", 
"01111001", 
"01111100", 
"01110100", 
"01100001", 
"01100110", 
"01101000", 
"01100110", 
"01110000", 
"10000011", 
"10001111", 
"10000001", 
"01101001", 
"01110111", 
"01110001", 
"01111100", 
"01110111", 
"01110111", 
"01110011", 
"01110110", 
"01011001", 
"01101011", 
"01101101", 
"10010000", 
"10000101", 
"10001011", 
"01111101", 
"01111111", 
"01011000", 
"01100110", 
"10000010", 
"10001010", 
"01101000", 
"01110110", 
"01101011", 
"01101000", 
"01110110", 
"10001010", 
"01111111", 
"01111010", 
"01110011", 
"01110101", 
"10001001", 
"01110111", 
"01110001", 
"10000011", 
"01111000", 
"10000000", 
"01100101", 
"01101110", 
"01101101", 
"01110011", 
"01110011", 
"01001010", 
"10010111", 
"01111010", 
"01010001", 
"10000001", 
"01111011", 
"01110111", 
"01100011", 
"10001101", 
"01111011", 
"10001111", 
"01100000", 
"01111101", 
"01110100", 
"10001010", 
"01111101", 
"10000111", 
"10001100", 
"10010111", 
"10001000", 
"01101000", 
"10010000", 
"01100011", 
"01101001", 
"01101011", 
"01111100", 
"10001100", 
"01110000", 
"01100001", 
"01111011", 
"10001110", 
"01111001", 
"01101010", 
"01100100", 
"01100110", 
"01101000", 
"01111111", 
"01111101", 
"01101011", 
"01101001", 
"01110110", 
"10001011", 
"01111110", 
"01100110", 
"01101110", 
"01111010", 
"10010010", 
"01101011", 
"10010001", 
"01010010", 
"01101100", 
"01101110", 
"01101010", 
"01110111", 
"01110000", 
"01001111", 
"01100100", 
"01101100", 
"01111011", 
"01001110", 
"10000111", 
"01100111", 
"10000010", 
"01110111", 
"01101100", 
"01100110", 
"01111001", 
"01111101", 
"10001100", 
"10000011", 
"10000100", 
"01110100", 
"01101101", 
"10001010", 
"10001101", 
"01110111", 
"01101000", 
"01101111", 
"10001010", 
"01111010", 
"10010001", 
"01101110", 
"01110001", 
"01100011", 
"01101011", 
"01110001", 
"01101001", 
"01111101", 
"01101001", 
"10010111", 
"01110010", 
"01110101", 
"10000000", 
"01110111", 
"10000010", 
"01100101", 
"01111011", 
"01101100", 
"01110010", 
"01110000", 
"01100110", 
"10001110", 
"01100011", 
"10001110", 
"01101010", 
"10001110", 
"10000011", 
"01111111", 
"10010000", 
"01111001", 
"10000011", 
"01110100", 
"01100100", 
"10000001", 
"01110010", 
"10000100", 
"01110001", 
"10010110", 
"01111000", 
"01011011", 
"01110000", 
"01111011", 
"01111011", 
"01000111", 
"01110111", 
"01101000", 
"01101011", 
"10001100", 
"01011011", 
"01110011", 
"01100111", 
"01111111", 
"10001110", 
"01110000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_107 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_107(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
