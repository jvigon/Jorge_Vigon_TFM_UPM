use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_9_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_9_LAYER;

architecture Behavioral of ROM_FC_84_9_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_9: ROM_ARRAY_PESOS_FC_84 := (
"10010001", 
"01100101", 
"10101010", 
"01101101", 
"01101010", 
"01111001", 
"01100101", 
"10000111", 
"10100100", 
"11000101", 
"01110000", 
"01111000", 
"01111110", 
"01100000", 
"10100010", 
"10001010", 
"01100010", 
"01111001", 
"01010111", 
"01110000", 
"10000110", 
"10000101", 
"01101001", 
"01110101", 
"01101111", 
"10010111", 
"01101110", 
"01110100", 
"01000001", 
"10011101", 
"10100101", 
"01111001", 
"01101000", 
"10011000", 
"01011110", 
"10100011", 
"01110110", 
"01100011", 
"01101100", 
"01111000", 
"10010011", 
"01101001", 
"01001000", 
"01100010", 
"10001110", 
"10010110", 
"01101010", 
"10000101", 
"01000111", 
"10001011", 
"01100111", 
"10011000", 
"10011111", 
"01110000", 
"10010011", 
"01110001", 
"10010000", 
"01111100", 
"01010101", 
"01110101", 
"01110101", 
"10010101", 
"01100001", 
"01011001", 
"10110000", 
"10000110", 
"10001001", 
"01111101", 
"01101011", 
"01011101", 
"01010010", 
"01010101", 
"10100100", 
"10000100", 
"01111111", 
"10010010", 
"01100100", 
"10001101", 
"10011000", 
"10000011", 
"01000011", 
"10001000", 
"01101010", 
"10001011", 
"10000111", 
"01011101", 
"10001010", 
"01101100", 
"10011100", 
"00111100", 
"01111101", 
"01101011", 
"10010111", 
"10000110", 
"01010000", 
"10000101", 
"10001010", 
"10010000", 
"10111111", 
"10001001", 
"01100011", 
"10001100", 
"10010000", 
"01010110", 
"10001110", 
"01110110", 
"10000110", 
"10001101", 
"01010110", 
"01110011", 
"01111110", 
"10000110", 
"01110100", 
"01001110", 
"10001000", 
"01100100", 
"10011011", 
"10110011", 
"01111001", 
"01101110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_9 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_9(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
