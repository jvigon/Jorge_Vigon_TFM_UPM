use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_60_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_60_LAYER;

architecture Behavioral of ROM_FC_120_60_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_60: ROM_ARRAY_PESOS_FC_120 := (
"10001100", 
"10111100", 
"01101011", 
"10000110", 
"01100001", 
"11011101", 
"01110110", 
"10010100", 
"01110100", 
"00111111", 
"01110111", 
"00010001", 
"01000001", 
"10101010", 
"10001000", 
"01101101", 
"10010111", 
"01101101", 
"01001000", 
"01101101", 
"01100111", 
"10100101", 
"10101000", 
"10010110", 
"10010101", 
"01100010", 
"01011100", 
"01000011", 
"01100010", 
"10010100", 
"01111100", 
"10000000", 
"10100010", 
"01000110", 
"01101010", 
"10001000", 
"01101001", 
"01110011", 
"10001110", 
"10001110", 
"01111001", 
"01110111", 
"01111011", 
"01010001", 
"01010010", 
"01001001", 
"01111101", 
"10001001", 
"10001110", 
"01000101", 
"10011001", 
"10001100", 
"10001101", 
"01110101", 
"10001001", 
"10100011", 
"10010000", 
"10010101", 
"01011000", 
"10000001", 
"10011100", 
"01110010", 
"01110110", 
"10001011", 
"10000000", 
"01101101", 
"10001011", 
"10011000", 
"01111001", 
"10001000", 
"01110001", 
"10000000", 
"10000000", 
"10000001", 
"01110101", 
"01011111", 
"10000001", 
"01011000", 
"01101000", 
"01111110", 
"10001010", 
"01100110", 
"10010001", 
"01111111", 
"10100110", 
"10001001", 
"01111100", 
"10010000", 
"10010000", 
"10010100", 
"01100101", 
"01010101", 
"10001101", 
"10000101", 
"01110011", 
"10010001", 
"01101110", 
"01010101", 
"10001101", 
"10000010", 
"10000101", 
"01111111", 
"10000100", 
"10000010", 
"01110011", 
"10010110", 
"01111000", 
"01011000", 
"01100000", 
"01001111", 
"01111011", 
"01111110", 
"01011010", 
"01110101", 
"01101011", 
"00010010", 
"10010101", 
"10000110", 
"01100011", 
"01011001", 
"01111001", 
"11001000", 
"01101010", 
"10100000", 
"10001010", 
"10000000", 
"10010010", 
"01110101", 
"01101010", 
"01011011", 
"01010000", 
"10010000", 
"10000111", 
"01111111", 
"01001101", 
"01011111", 
"10000001", 
"10010000", 
"01100101", 
"01000011", 
"01100100", 
"01110101", 
"01111011", 
"10001011", 
"01111100", 
"01111111", 
"10001000", 
"01100111", 
"01110000", 
"01011110", 
"01101100", 
"01110111", 
"10011010", 
"10000000", 
"10000110", 
"01011100", 
"10011011", 
"01111101", 
"01111111", 
"01101100", 
"01100100", 
"10011110", 
"01101100", 
"01000100", 
"01111111", 
"01111111", 
"01010100", 
"01010100", 
"10000000", 
"01101111", 
"01100010", 
"01110101", 
"10001110", 
"10101000", 
"10000111", 
"01110100", 
"01110110", 
"10100010", 
"10000111", 
"00110100", 
"10010100", 
"10010100", 
"10010001", 
"01101101", 
"01110000", 
"01101100", 
"10001010", 
"10010100", 
"10011110", 
"10100001", 
"01111100", 
"01110101", 
"10000111", 
"10001010", 
"01101101", 
"01001101", 
"01110011", 
"10000001", 
"01000110", 
"01110001", 
"01100111", 
"10011000", 
"01010100", 
"01101110", 
"10000110", 
"10010101", 
"01110011", 
"10000010", 
"01111011", 
"10011010", 
"01011111", 
"01101101", 
"10000011", 
"01011100", 
"01011110", 
"01101100", 
"10000001", 
"10001001", 
"10010000", 
"10010100", 
"10000100", 
"10000010", 
"01110101", 
"10001110", 
"01110011", 
"01111010", 
"01110010", 
"01010111", 
"01101100", 
"10001100", 
"01111101", 
"10000010", 
"10010111", 
"10000111", 
"01000011", 
"01100010", 
"01111100", 
"01111101", 
"01101101", 
"10010011", 
"01000110", 
"01111010", 
"01101100", 
"01011011", 
"01110100", 
"01110010", 
"01101101", 
"10000101", 
"01100110", 
"01011000", 
"01100100", 
"01010101", 
"10111100", 
"10000010", 
"10001010", 
"01101011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_60: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_60(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
