use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_87_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_87_LAYER;

architecture Behavioral of ROM_FC_120_87_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_87: ROM_ARRAY_PESOS_FC_120 := (
"10111101", 
"01101111", 
"01110110", 
"01101111", 
"01111101", 
"10101100", 
"01011010", 
"10000111", 
"01100010", 
"01111011", 
"01111101", 
"01011000", 
"01011101", 
"01111100", 
"01111101", 
"10000101", 
"10001000", 
"01111110", 
"10011101", 
"01100101", 
"10101101", 
"01011110", 
"10000101", 
"10001100", 
"10001010", 
"01111111", 
"01111001", 
"01110010", 
"01110000", 
"10111101", 
"01110011", 
"01111101", 
"01001010", 
"01110101", 
"10000101", 
"01001111", 
"11111111", 
"01000100", 
"10001101", 
"01010010", 
"01111000", 
"01111001", 
"01000010", 
"10011000", 
"10010001", 
"01110000", 
"10000100", 
"01111000", 
"10010001", 
"10100010", 
"10010011", 
"01111011", 
"01101101", 
"01111000", 
"10100010", 
"01110101", 
"10001100", 
"01100100", 
"10001101", 
"01111001", 
"01110101", 
"10000001", 
"10101011", 
"10000011", 
"01010100", 
"01111001", 
"00101100", 
"00100111", 
"11000010", 
"01101110", 
"01101001", 
"01111100", 
"01010000", 
"01111111", 
"01111110", 
"01110110", 
"10001110", 
"10001110", 
"01110010", 
"10010111", 
"00100111", 
"01110110", 
"01101111", 
"01101101", 
"10010111", 
"01110101", 
"01111111", 
"10011111", 
"01011110", 
"01101101", 
"01100101", 
"10011100", 
"10001000", 
"10011001", 
"10001110", 
"01110100", 
"01110001", 
"10000100", 
"10010000", 
"01101100", 
"10100010", 
"01010111", 
"01101101", 
"01110100", 
"01101001", 
"01110011", 
"01000010", 
"01111100", 
"10111001", 
"01010000", 
"01101001", 
"01110011", 
"10000110", 
"10100111", 
"01101010", 
"01011100", 
"10100100", 
"01111000", 
"00101100", 
"10011011", 
"01110011", 
"10101101", 
"01001010", 
"01101101", 
"01110100", 
"01100111", 
"10000010", 
"01111101", 
"01100001", 
"01110000", 
"10011101", 
"01111011", 
"01100101", 
"01100100", 
"01000101", 
"01001010", 
"10001111", 
"01011000", 
"01101111", 
"10000101", 
"01110001", 
"11000000", 
"10000010", 
"01111000", 
"01000100", 
"01011110", 
"10000101", 
"01100010", 
"11001001", 
"01101110", 
"01101010", 
"01101001", 
"10101010", 
"01001100", 
"01000101", 
"01010111", 
"10100101", 
"01011110", 
"10100000", 
"10000001", 
"01011011", 
"01011011", 
"10000010", 
"10010001", 
"10010110", 
"10001110", 
"01100111", 
"10000100", 
"01011100", 
"01101010", 
"10100110", 
"01001001", 
"01111100", 
"11011001", 
"01100100", 
"10000111", 
"01111001", 
"01001000", 
"01100100", 
"10010011", 
"10000010", 
"10000100", 
"01010101", 
"10110101", 
"01011000", 
"10000101", 
"00110011", 
"01011010", 
"01100111", 
"01100011", 
"10000100", 
"10000010", 
"01011100", 
"10000110", 
"10000010", 
"10011011", 
"10100100", 
"01010100", 
"01111001", 
"01000011", 
"01111111", 
"10000011", 
"10001001", 
"01110100", 
"10011000", 
"11111111", 
"01100001", 
"01110001", 
"00100111", 
"10011110", 
"01110111", 
"10001011", 
"10000010", 
"01011001", 
"10111010", 
"01100011", 
"01101001", 
"01110110", 
"00100110", 
"01110011", 
"11000011", 
"01111001", 
"01101110", 
"10001010", 
"01110101", 
"10010010", 
"10000010", 
"10001110", 
"10000101", 
"01110101", 
"01100111", 
"10011010", 
"01000000", 
"00110110", 
"01111000", 
"01111011", 
"01101111", 
"10010010", 
"01111111", 
"01110001", 
"10010001", 
"10101010", 
"01000010", 
"01001100", 
"10000100", 
"01111111", 
"10000110", 
"01111101", 
"10011100", 
"00101100", 
"01111011", 
"01100010", 
"01101000", 
"11001100", 
"01101011", 
"01111000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_87: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_87(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
