use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_106_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_106_LAYER;

architecture Behavioral of ROM_FC_120_106_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_106: ROM_ARRAY_PESOS_FC_120 := (
"01101110", 
"01111101", 
"01100101", 
"10000111", 
"01110111", 
"01111111", 
"01101100", 
"01100000", 
"10000011", 
"01101111", 
"10000000", 
"01111110", 
"01010101", 
"01110110", 
"10000011", 
"10001111", 
"01101011", 
"01100110", 
"01111111", 
"10010110", 
"10000000", 
"01010100", 
"01101001", 
"01110111", 
"01110111", 
"01101011", 
"01011101", 
"10000011", 
"01100111", 
"10101000", 
"01111000", 
"01111011", 
"01100010", 
"01100000", 
"10001100", 
"01111001", 
"01101111", 
"01110101", 
"01110111", 
"01011010", 
"10001110", 
"10000110", 
"10001111", 
"01110111", 
"01111101", 
"01101001", 
"01101011", 
"10001111", 
"01110011", 
"01101111", 
"10000110", 
"01011111", 
"01111011", 
"01101000", 
"01011100", 
"01011110", 
"01101111", 
"01110100", 
"01101010", 
"01111100", 
"10000110", 
"01111011", 
"10001010", 
"01111000", 
"01100100", 
"01110101", 
"01101000", 
"10001110", 
"01111111", 
"10000001", 
"01111101", 
"01111110", 
"01110011", 
"01011001", 
"01110001", 
"01011010", 
"01111011", 
"10000100", 
"10000111", 
"10001000", 
"01101111", 
"01111011", 
"01101010", 
"01011111", 
"01111010", 
"10001000", 
"10000011", 
"01110001", 
"10000000", 
"01100010", 
"01001110", 
"01101101", 
"01101000", 
"01001111", 
"10001001", 
"10000001", 
"01001000", 
"01110110", 
"01111100", 
"01111001", 
"01101010", 
"01110010", 
"01111110", 
"01101011", 
"10000100", 
"01110111", 
"01100101", 
"01101011", 
"01100100", 
"10101010", 
"10000000", 
"01110100", 
"01100011", 
"01110010", 
"01111100", 
"01100011", 
"01111000", 
"01111010", 
"10000101", 
"01101010", 
"10000101", 
"10000000", 
"01100001", 
"10000111", 
"10010110", 
"01101010", 
"01101101", 
"01111100", 
"01101011", 
"10010011", 
"10001001", 
"01111000", 
"10001000", 
"01111010", 
"01110001", 
"01111110", 
"01101011", 
"01011111", 
"10001000", 
"01101100", 
"10010011", 
"01011010", 
"01111010", 
"10001001", 
"10001011", 
"10000111", 
"01110011", 
"01111011", 
"10001010", 
"10000110", 
"01101111", 
"01111000", 
"10001110", 
"10000111", 
"01101001", 
"01111000", 
"10011000", 
"01100111", 
"01110001", 
"10000010", 
"01111101", 
"01111110", 
"10000010", 
"10001100", 
"10000111", 
"01110111", 
"10000110", 
"01100001", 
"10001001", 
"10000111", 
"01110011", 
"01111110", 
"01111011", 
"10011010", 
"10001010", 
"01100101", 
"10000101", 
"01110101", 
"01011111", 
"01110101", 
"01111001", 
"01011111", 
"10001110", 
"01111111", 
"01111101", 
"01111101", 
"01010110", 
"01111101", 
"01100111", 
"10001100", 
"10001101", 
"01111011", 
"01111010", 
"10001011", 
"01001011", 
"01101110", 
"01101111", 
"01101001", 
"10001101", 
"10000000", 
"01111111", 
"10000000", 
"01100111", 
"01101101", 
"01011111", 
"01100100", 
"01110100", 
"10001011", 
"01111011", 
"01101101", 
"01001110", 
"01011000", 
"01101110", 
"10000010", 
"10010100", 
"10000110", 
"10010100", 
"01110010", 
"01111000", 
"01100110", 
"01100101", 
"01001010", 
"10000100", 
"01110110", 
"01110110", 
"01100010", 
"01110110", 
"10001100", 
"10010010", 
"01100011", 
"01111101", 
"01101110", 
"01110111", 
"01010101", 
"10001100", 
"01100000", 
"01101011", 
"01111100", 
"10010010", 
"10000000", 
"01011001", 
"01101111", 
"10001000", 
"10011100", 
"01110011", 
"01001101", 
"10001000", 
"01100100", 
"01111010", 
"01101111", 
"01100110", 
"01101010", 
"01001110", 
"10010101", 
"01111111", 
"01111011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_106 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_106(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
