use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_47_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_47_LAYER;

architecture Behavioral of ROM_FC_84_47_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_47: ROM_ARRAY_PESOS_FC_84 := (
"10000010", 
"01010011", 
"10001111", 
"01110100", 
"01011000", 
"10001110", 
"01100000", 
"10011010", 
"01101111", 
"10001000", 
"10000011", 
"01110101", 
"10000010", 
"01110011", 
"10001110", 
"10001001", 
"10001110", 
"10001110", 
"01011000", 
"01000000", 
"01101100", 
"01101000", 
"10100000", 
"01101000", 
"10001101", 
"10010111", 
"10100000", 
"01110100", 
"01100000", 
"10000100", 
"10010010", 
"01001100", 
"01101110", 
"10000111", 
"10110010", 
"01110010", 
"11000001", 
"10100101", 
"01011000", 
"01001000", 
"10010100", 
"10001001", 
"10000110", 
"01001010", 
"10101010", 
"01010000", 
"01110101", 
"01111001", 
"01110100", 
"10001010", 
"01101000", 
"10111010", 
"01101001", 
"10000011", 
"01111110", 
"10100101", 
"01110011", 
"01110100", 
"01101111", 
"00111101", 
"10000100", 
"10010001", 
"10001100", 
"10011011", 
"01110110", 
"10000101", 
"01111101", 
"10010101", 
"10000000", 
"01011000", 
"01100001", 
"01010101", 
"00110110", 
"01101111", 
"01111111", 
"01110110", 
"10100010", 
"01111101", 
"10011001", 
"10011011", 
"10110000", 
"10000001", 
"01110001", 
"01010100", 
"10100000", 
"01100001", 
"01010000", 
"10101111", 
"01111101", 
"00101111", 
"10111110", 
"01111011", 
"01110010", 
"00111110", 
"10110111", 
"10100111", 
"10000100", 
"10010101", 
"10000001", 
"10101001", 
"10010100", 
"10000010", 
"10101100", 
"10001000", 
"01100010", 
"10000110", 
"10100011", 
"01101110", 
"01001000", 
"01010011", 
"10100110", 
"01100111", 
"01111111", 
"10100001", 
"10000111", 
"00111101", 
"01110111", 
"01010001", 
"10000001", 
"10000011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_47: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_47(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
