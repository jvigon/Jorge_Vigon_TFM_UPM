use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_43_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_43_LAYER;

architecture Behavioral of ROM_FC_120_43_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_43: ROM_ARRAY_PESOS_FC_120 := (
"01110101", 
"10000011", 
"10110110", 
"10111100", 
"01011111", 
"01110110", 
"01010101", 
"01011111", 
"10001110", 
"10101011", 
"01110010", 
"10100011", 
"10000101", 
"11010001", 
"10010001", 
"10010000", 
"10011001", 
"10111000", 
"01101110", 
"01101100", 
"01110011", 
"01010101", 
"00110101", 
"10011011", 
"01110110", 
"10011010", 
"10010000", 
"10010000", 
"10001111", 
"11000111", 
"01110111", 
"10011001", 
"10101101", 
"10000001", 
"01100010", 
"01101001", 
"01111000", 
"10011110", 
"01000011", 
"10000001", 
"10000101", 
"10011111", 
"01010001", 
"01101011", 
"10010101", 
"10001011", 
"01110011", 
"01110101", 
"10010011", 
"10001000", 
"10011100", 
"01011100", 
"01111000", 
"10100100", 
"10011010", 
"10101101", 
"01110010", 
"01101001", 
"01100010", 
"01000010", 
"10101111", 
"01101100", 
"10001011", 
"10000011", 
"10000101", 
"11001100", 
"10001010", 
"00010010", 
"01011101", 
"10100010", 
"01001010", 
"01110101", 
"10001001", 
"10100001", 
"10110110", 
"10110011", 
"10010000", 
"01000001", 
"01111110", 
"10000111", 
"01101110", 
"10100111", 
"01011110", 
"00001010", 
"01101111", 
"01111001", 
"01101001", 
"01110110", 
"01101101", 
"10011001", 
"10110000", 
"10101000", 
"10000001", 
"10111010", 
"01110100", 
"01110010", 
"01111000", 
"10001000", 
"01100001", 
"01100110", 
"10001101", 
"01110000", 
"10001100", 
"01010111", 
"10001001", 
"10101001", 
"01101010", 
"10011100", 
"10010100", 
"10010010", 
"01101111", 
"10000111", 
"10011001", 
"10001101", 
"10000110", 
"10010001", 
"01101111", 
"01100111", 
"00111010", 
"01111010", 
"10000111", 
"10010110", 
"10010110", 
"01100001", 
"10011010", 
"01100110", 
"01101011", 
"10010000", 
"10000101", 
"01111101", 
"01010000", 
"00100001", 
"01101101", 
"10101010", 
"01100111", 
"10111110", 
"01111101", 
"01001110", 
"10011110", 
"10001101", 
"10010101", 
"10011011", 
"01101100", 
"01111001", 
"10010110", 
"01101100", 
"10001001", 
"01000101", 
"10000111", 
"10000101", 
"01110100", 
"10011110", 
"10001110", 
"10000100", 
"01100101", 
"01110001", 
"10000110", 
"10100101", 
"10000101", 
"10000010", 
"10001110", 
"01111010", 
"10001010", 
"01111100", 
"01101110", 
"10001110", 
"10011111", 
"01110101", 
"10011001", 
"10010101", 
"01101101", 
"11001011", 
"01110011", 
"01000110", 
"01100111", 
"01110100", 
"10011001", 
"01101110", 
"10110000", 
"10000111", 
"10001011", 
"01111101", 
"10000000", 
"01110101", 
"01111101", 
"10000001", 
"01110111", 
"10100101", 
"10011111", 
"01111111", 
"01111100", 
"01111000", 
"01101100", 
"01110010", 
"00101010", 
"00100000", 
"01110010", 
"10010101", 
"10101101", 
"10010010", 
"10010001", 
"01100000", 
"01110111", 
"01111101", 
"01000111", 
"10011101", 
"10001010", 
"01100111", 
"10101010", 
"01100000", 
"00101110", 
"00011100", 
"01111001", 
"10001011", 
"10000010", 
"01111000", 
"01111001", 
"01011001", 
"10010101", 
"10001011", 
"01010100", 
"01111110", 
"01111011", 
"01111011", 
"01100110", 
"01100010", 
"01010111", 
"00111000", 
"01111111", 
"10001100", 
"10101010", 
"10001111", 
"10010111", 
"01101101", 
"10100000", 
"01100011", 
"10100100", 
"01100111", 
"01110000", 
"01101001", 
"01101000", 
"01011110", 
"01110010", 
"01100000", 
"01110011", 
"01110001", 
"10000010", 
"01111111", 
"10000110", 
"01101001", 
"10111011", 
"01000010", 
"01011000", 
"01101101", 
"10000011", 
"01100011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_43: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_43(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
