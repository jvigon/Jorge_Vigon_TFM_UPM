use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_93_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_93_LAYER;

architecture Behavioral of ROM_FC_120_93_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_93: ROM_ARRAY_PESOS_FC_120 := (
"01110101", 
"10100110", 
"00100111", 
"01011001", 
"10000101", 
"10100101", 
"10001110", 
"11000000", 
"10000010", 
"01011110", 
"01110111", 
"01011100", 
"01000111", 
"00111000", 
"01101110", 
"01111110", 
"10101010", 
"01111000", 
"01100101", 
"01001101", 
"01010111", 
"10000001", 
"10100011", 
"11011001", 
"01101101", 
"01111111", 
"10000110", 
"00011111", 
"01011000", 
"01010111", 
"01111100", 
"10011000", 
"10111101", 
"10011111", 
"01110111", 
"01101000", 
"10000010", 
"01111101", 
"10101000", 
"10011110", 
"01110001", 
"01101010", 
"01101101", 
"01111010", 
"10000000", 
"01011100", 
"01101101", 
"10001000", 
"10010010", 
"01110101", 
"01100001", 
"10000000", 
"10000001", 
"10000100", 
"01100110", 
"10110110", 
"10000010", 
"01100010", 
"01111000", 
"01101001", 
"10001100", 
"10000000", 
"01101100", 
"10001101", 
"10001010", 
"01010000", 
"01100000", 
"01101011", 
"01100100", 
"10011110", 
"01111101", 
"10010111", 
"10011100", 
"01011000", 
"01110011", 
"00000000", 
"01101111", 
"00001000", 
"10000111", 
"01101011", 
"11000000", 
"01001010", 
"10001010", 
"01110100", 
"10001011", 
"10001000", 
"01111001", 
"10001001", 
"01010000", 
"01110010", 
"10010011", 
"01010100", 
"01101111", 
"01101111", 
"10000001", 
"01110110", 
"10011111", 
"10100111", 
"01100111", 
"10000000", 
"10111110", 
"01000011", 
"10010000", 
"10001001", 
"01110100", 
"10010111", 
"01110111", 
"10100011", 
"01110010", 
"10011000", 
"01110110", 
"10000000", 
"00010110", 
"11000000", 
"01111101", 
"01101000", 
"10101101", 
"01100000", 
"01111011", 
"01101110", 
"10000110", 
"00101111", 
"01100001", 
"10001010", 
"10110011", 
"10101110", 
"10000111", 
"10000001", 
"01010001", 
"10000000", 
"01110011", 
"10001010", 
"01101010", 
"10100101", 
"01101100", 
"01111001", 
"01110010", 
"00100011", 
"10010100", 
"00100110", 
"00100010", 
"01011010", 
"01111101", 
"10000000", 
"01110111", 
"00111100", 
"01111101", 
"10010100", 
"10010101", 
"01101110", 
"10011111", 
"01110111", 
"01100010", 
"01010111", 
"10110011", 
"01010010", 
"01111000", 
"10010001", 
"10000111", 
"10000010", 
"01010101", 
"01010111", 
"10011010", 
"10010110", 
"10010101", 
"01100011", 
"01101000", 
"00110111", 
"10000110", 
"01100101", 
"01110110", 
"01011101", 
"10011001", 
"01110110", 
"01110100", 
"10010001", 
"10101010", 
"10110111", 
"10010111", 
"01001101", 
"10001110", 
"01100101", 
"10000000", 
"01001110", 
"10010111", 
"01110101", 
"01101001", 
"01101000", 
"11010110", 
"10100011", 
"10000110", 
"10000010", 
"10001100", 
"01111000", 
"10010011", 
"10001111", 
"01011111", 
"10101100", 
"01100001", 
"01010000", 
"10001000", 
"01011101", 
"01110110", 
"00110011", 
"00100100", 
"10100100", 
"10000110", 
"01111001", 
"00110011", 
"01010010", 
"10110101", 
"10100101", 
"10000011", 
"01010101", 
"10010011", 
"01100001", 
"10001101", 
"10010000", 
"10100001", 
"00100011", 
"01110101", 
"10101010", 
"10000101", 
"01110101", 
"01101011", 
"01110101", 
"10011010", 
"10101011", 
"01011100", 
"10100011", 
"10000110", 
"10100100", 
"01110011", 
"10011010", 
"10010001", 
"01101110", 
"10000110", 
"10011100", 
"01110110", 
"01111010", 
"01111011", 
"10001100", 
"01111011", 
"10101011", 
"01111101", 
"10001010", 
"10101010", 
"10100100", 
"10001110", 
"10001111", 
"01011101", 
"01100001", 
"01110011", 
"01011000", 
"01110110", 
"01111000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_93: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_93(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
