use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_25_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_25_LAYER;

architecture Behavioral of ROM_FC_120_25_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_25: ROM_ARRAY_PESOS_FC_120 := (
"10011100", 
"00110111", 
"01110010", 
"01111010", 
"01111110", 
"10101001", 
"01101000", 
"01100011", 
"01101001", 
"10000110", 
"10011111", 
"01010110", 
"01100000", 
"01111000", 
"01110111", 
"10001000", 
"01101110", 
"01001010", 
"01001010", 
"10001000", 
"10001001", 
"01101011", 
"01111110", 
"10101001", 
"01110110", 
"01110000", 
"01110110", 
"01111111", 
"00101001", 
"10101010", 
"10001111", 
"01110100", 
"01011010", 
"01111011", 
"01011001", 
"01110011", 
"01101001", 
"00111110", 
"10000010", 
"01001001", 
"01110010", 
"01101101", 
"01010001", 
"10011001", 
"01001011", 
"01100110", 
"01110110", 
"10000010", 
"01111100", 
"01110101", 
"10001111", 
"01111101", 
"10000001", 
"01100100", 
"10001101", 
"01110111", 
"10000110", 
"10001000", 
"01111000", 
"10000111", 
"10001111", 
"00110000", 
"10000100", 
"01110001", 
"10000110", 
"00111000", 
"00111000", 
"10111111", 
"01110000", 
"10011101", 
"01011100", 
"10010001", 
"10011111", 
"01000010", 
"10100010", 
"01111011", 
"01010001", 
"01110011", 
"10000110", 
"01111110", 
"01000101", 
"00110000", 
"01100101", 
"01101011", 
"10000111", 
"01101110", 
"10000100", 
"10001110", 
"01100110", 
"01011111", 
"01000000", 
"01101111", 
"01111010", 
"01111011", 
"01101011", 
"01110001", 
"01100010", 
"10001000", 
"01110101", 
"01101111", 
"10000011", 
"00110011", 
"01101001", 
"01110111", 
"01101010", 
"01111001", 
"00111101", 
"01101010", 
"10010010", 
"01110001", 
"01111011", 
"10001100", 
"01001001", 
"10001100", 
"01100100", 
"10000110", 
"10001000", 
"01100111", 
"10010001", 
"01111101", 
"10001111", 
"01101001", 
"01100110", 
"10010111", 
"01100100", 
"01011010", 
"01110110", 
"01111001", 
"01000110", 
"01001100", 
"01100010", 
"10010101", 
"01110110", 
"11001000", 
"01110001", 
"01000011", 
"01111100", 
"10001001", 
"10101101", 
"01000101", 
"01001110", 
"01011001", 
"10001111", 
"10000100", 
"01101100", 
"01111011", 
"10001110", 
"01111010", 
"01101101", 
"01010011", 
"00111001", 
"01101011", 
"01110010", 
"10000010", 
"01100010", 
"00101111", 
"01110111", 
"10011000", 
"01111100", 
"10000110", 
"01000111", 
"01110110", 
"01011010", 
"01111011", 
"10001100", 
"01110100", 
"10010100", 
"10011010", 
"10000001", 
"10000100", 
"01011111", 
"10001001", 
"01010011", 
"01100110", 
"10001010", 
"01110001", 
"01001101", 
"01110010", 
"01110001", 
"10010101", 
"01111010", 
"01011101", 
"10100110", 
"01001000", 
"10000111", 
"01111000", 
"01100011", 
"10101101", 
"10001110", 
"01110110", 
"01111101", 
"10000011", 
"01011100", 
"01111101", 
"01100000", 
"01001111", 
"01100110", 
"01110001", 
"01100001", 
"01100011", 
"01111111", 
"01001100", 
"01001101", 
"01011110", 
"01111010", 
"10010000", 
"10000001", 
"01111010", 
"01011001", 
"01100100", 
"10000000", 
"10010110", 
"01110010", 
"01101000", 
"01010110", 
"01011100", 
"01101100", 
"01010100", 
"01111001", 
"01110010", 
"10000011", 
"10001000", 
"10000000", 
"01111110", 
"10000000", 
"01011101", 
"01101111", 
"10000100", 
"10000010", 
"01001110", 
"10010010", 
"01010100", 
"10000011", 
"01101001", 
"10000001", 
"10001110", 
"10100001", 
"01010110", 
"10000011", 
"01111011", 
"10000100", 
"01001010", 
"01111001", 
"10001010", 
"01101101", 
"01110001", 
"10011110", 
"01111101", 
"10001101", 
"10001100", 
"01001110", 
"01011100", 
"01010100", 
"10000000", 
"10001000", 
"01111110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_25: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_25(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
