use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_53_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_53_LAYER;

architecture Behavioral of ROM_FC_120_53_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_53: ROM_ARRAY_PESOS_FC_120 := (
"01111010", 
"01101110", 
"01111111", 
"10000100", 
"01100101", 
"01001011", 
"10010110", 
"10000011", 
"10001110", 
"10011011", 
"01110010", 
"00100110", 
"01111000", 
"10010010", 
"10001011", 
"10000001", 
"01111000", 
"10000001", 
"10001010", 
"00101010", 
"01111111", 
"01100101", 
"01101100", 
"01110100", 
"10001000", 
"10011100", 
"10100001", 
"01101101", 
"01100101", 
"10011101", 
"01111000", 
"01111110", 
"01110111", 
"01110011", 
"10000110", 
"10000010", 
"01111001", 
"01101001", 
"01100010", 
"10001001", 
"10001111", 
"01110011", 
"10010000", 
"10011010", 
"01110111", 
"10101000", 
"01111011", 
"10010111", 
"01101101", 
"01111101", 
"01101001", 
"10111101", 
"10010001", 
"01110100", 
"01111000", 
"01111011", 
"01111011", 
"00111101", 
"01110001", 
"01110111", 
"10101101", 
"10110101", 
"10011000", 
"10001110", 
"10000101", 
"10000110", 
"01111001", 
"01011100", 
"10000101", 
"10010110", 
"01101001", 
"01110101", 
"10000110", 
"01111011", 
"10110111", 
"01001111", 
"10000100", 
"01110000", 
"10001111", 
"10001110", 
"10010100", 
"01111011", 
"01110000", 
"01101000", 
"01111100", 
"01011001", 
"01001101", 
"01110100", 
"01110011", 
"01111001", 
"01110111", 
"01010110", 
"10000011", 
"10000111", 
"10000011", 
"10000101", 
"01110000", 
"01111001", 
"01110111", 
"01011001", 
"01110101", 
"01101111", 
"01100111", 
"01100111", 
"10010000", 
"01110011", 
"01100011", 
"10101010", 
"01100001", 
"10001010", 
"10010000", 
"01111011", 
"01101111", 
"10000101", 
"01111001", 
"10101010", 
"10010001", 
"01110010", 
"10100000", 
"01110010", 
"10001001", 
"01110101", 
"01100010", 
"10110001", 
"10000100", 
"01110011", 
"01110110", 
"10100100", 
"10001010", 
"10001110", 
"10011110", 
"10011101", 
"10000100", 
"10110010", 
"01111000", 
"01111010", 
"10001100", 
"01000110", 
"10101110", 
"00001000", 
"01000000", 
"01111000", 
"01111010", 
"01111001", 
"10000111", 
"01101101", 
"01110000", 
"01111011", 
"10000110", 
"10001010", 
"01010101", 
"10001001", 
"10001111", 
"01110110", 
"01101011", 
"01001001", 
"01001011", 
"10101000", 
"01110011", 
"01110110", 
"01111000", 
"01111011", 
"01111010", 
"01101100", 
"01110111", 
"01111100", 
"10100010", 
"01111011", 
"01110111", 
"10010000", 
"01100111", 
"10011101", 
"10001110", 
"01101111", 
"10010010", 
"01101100", 
"01101000", 
"10001100", 
"10010010", 
"01001110", 
"10000000", 
"01110001", 
"10010101", 
"01100010", 
"01101111", 
"10001010", 
"01110000", 
"10000111", 
"10000101", 
"01010100", 
"01111010", 
"01110110", 
"01111011", 
"10100111", 
"01111100", 
"10011100", 
"01110110", 
"10010100", 
"01010110", 
"01100011", 
"01111101", 
"01001111", 
"10010001", 
"01001010", 
"01110011", 
"10000110", 
"10001100", 
"01111000", 
"10001100", 
"10000101", 
"01101000", 
"01100001", 
"10001010", 
"01110010", 
"10010011", 
"01101011", 
"01110001", 
"01101010", 
"10001010", 
"01011101", 
"01100110", 
"10010110", 
"01111110", 
"01111101", 
"01110011", 
"01101011", 
"01101101", 
"01111011", 
"01110100", 
"01101001", 
"10001101", 
"01101100", 
"10000011", 
"01111100", 
"01110101", 
"10010100", 
"10110110", 
"01110010", 
"01110100", 
"01100110", 
"10010110", 
"10001110", 
"10000010", 
"00100110", 
"10010101", 
"01100000", 
"10001110", 
"01111110", 
"10001101", 
"10001110", 
"01111000", 
"10010001", 
"10011100", 
"01111001", 
"01110100", 
"01110000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_53: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_53(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
