use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_59_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_59_LAYER;

architecture Behavioral of ROM_FC_84_59_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_59: ROM_ARRAY_PESOS_FC_84 := (
"01110010", 
"01001101", 
"01010001", 
"10001001", 
"01101111", 
"10000001", 
"01110100", 
"01000111", 
"10000110", 
"01111010", 
"10010101", 
"10010000", 
"01100010", 
"10001000", 
"00110010", 
"01110011", 
"10001110", 
"01110110", 
"01110001", 
"10100000", 
"01011111", 
"01101111", 
"10001000", 
"01111000", 
"10001110", 
"01011100", 
"01101010", 
"01111110", 
"10011101", 
"01111111", 
"10011010", 
"01011101", 
"10011001", 
"10010000", 
"10000011", 
"01000001", 
"01100011", 
"10100100", 
"01110110", 
"01100000", 
"01100010", 
"01101110", 
"01100001", 
"01100010", 
"01101100", 
"01111110", 
"01110100", 
"10010110", 
"01101101", 
"01101101", 
"01011110", 
"01110001", 
"10001101", 
"10001011", 
"01011111", 
"10111011", 
"10100100", 
"10000100", 
"01010101", 
"01110110", 
"01010000", 
"01001000", 
"01110110", 
"10100110", 
"01101000", 
"01110001", 
"01110100", 
"01111000", 
"01110010", 
"01101110", 
"01111100", 
"00111010", 
"00100111", 
"10010010", 
"01110001", 
"10010111", 
"01101000", 
"10000010", 
"01101101", 
"10000001", 
"01001110", 
"01110111", 
"10001011", 
"01010110", 
"01101011", 
"10001100", 
"01010000", 
"10101100", 
"10010000", 
"10001011", 
"10110100", 
"01101011", 
"01110100", 
"01101001", 
"01110101", 
"10011000", 
"01010111", 
"01101010", 
"10000111", 
"10011000", 
"01110111", 
"01111100", 
"10101101", 
"10000001", 
"01001010", 
"01100111", 
"10001101", 
"10011111", 
"01110001", 
"01101111", 
"10001100", 
"01111001", 
"10000110", 
"01011100", 
"01111000", 
"01011111", 
"10001000", 
"10101110", 
"10000010", 
"01111001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_59: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_59(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
