use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_17_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_17_LAYER;

architecture Behavioral of ROM_FC_84_17_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_17: ROM_ARRAY_PESOS_FC_84 := (
"10010000", 
"01111101", 
"10010101", 
"10000001", 
"01110001", 
"10001000", 
"10011001", 
"01111110", 
"10000110", 
"01100001", 
"01110001", 
"01010000", 
"01111011", 
"10001100", 
"01110101", 
"10011100", 
"01001000", 
"01111010", 
"10011010", 
"10101111", 
"10100000", 
"10101101", 
"10001010", 
"10000010", 
"10010000", 
"10000100", 
"01111001", 
"10000000", 
"01001100", 
"10010011", 
"10001000", 
"01000100", 
"10000001", 
"10000000", 
"01001100", 
"01110110", 
"01111101", 
"01111110", 
"01101011", 
"01011110", 
"01100100", 
"10001100", 
"01001110", 
"01010010", 
"01110101", 
"10101001", 
"01011110", 
"10010011", 
"01111000", 
"01111011", 
"10000111", 
"01100011", 
"01101011", 
"01010101", 
"10100101", 
"10001100", 
"01110100", 
"10001111", 
"10011110", 
"01110110", 
"10100000", 
"10010011", 
"10010101", 
"10011100", 
"10011111", 
"01101010", 
"01101110", 
"10010111", 
"01110110", 
"01011001", 
"01000111", 
"10110100", 
"10101111", 
"10010100", 
"10010010", 
"01101111", 
"01110011", 
"01110000", 
"01101111", 
"01001000", 
"10001000", 
"01100001", 
"01011101", 
"10011001", 
"10010001", 
"01100111", 
"01000000", 
"01110011", 
"10011101", 
"01010001", 
"10000001", 
"10001001", 
"10011011", 
"10110110", 
"01111000", 
"01110001", 
"01011001", 
"10000010", 
"10000100", 
"01110111", 
"10001001", 
"01101111", 
"01110011", 
"01010000", 
"01111000", 
"01110111", 
"01111000", 
"01101010", 
"10000101", 
"10110100", 
"11000111", 
"10001001", 
"10001010", 
"10100100", 
"01111001", 
"01000010", 
"10000100", 
"10100110", 
"01110101", 
"01111111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_17 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_17(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
