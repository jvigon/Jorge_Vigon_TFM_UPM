use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_51_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_51_LAYER;

architecture Behavioral of ROM_FC_120_51_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_51: ROM_ARRAY_PESOS_FC_120 := (
"10000100", 
"01010010", 
"01111000", 
"10010010", 
"10000010", 
"01101011", 
"10001110", 
"10000011", 
"01110101", 
"10010011", 
"01010010", 
"10000010", 
"10010111", 
"10100110", 
"10000010", 
"01111110", 
"10010001", 
"01011110", 
"01011010", 
"01010011", 
"01101001", 
"01100011", 
"01010001", 
"10000110", 
"01110110", 
"11000110", 
"01100011", 
"01101000", 
"01111011", 
"10000111", 
"10000111", 
"10001111", 
"01111111", 
"10000000", 
"01101111", 
"01101000", 
"01110001", 
"00111101", 
"01011011", 
"01100100", 
"01110011", 
"10111011", 
"01110001", 
"01111110", 
"01101100", 
"01101001", 
"01101110", 
"01111100", 
"01111010", 
"01101011", 
"01101100", 
"01011111", 
"10001010", 
"01011111", 
"10011001", 
"01100111", 
"10000100", 
"01100100", 
"01101101", 
"01010111", 
"10011111", 
"01011001", 
"10000110", 
"01110100", 
"10001110", 
"01101100", 
"01101111", 
"01101100", 
"10001001", 
"10001100", 
"01011011", 
"10001100", 
"01111101", 
"01111000", 
"01100000", 
"01111100", 
"01100010", 
"01100111", 
"10000111", 
"01111100", 
"10001101", 
"10000101", 
"01110111", 
"01000111", 
"01111100", 
"01100001", 
"01110011", 
"10001000", 
"01101101", 
"10010001", 
"01101001", 
"10001011", 
"10011011", 
"01010100", 
"01110000", 
"01111111", 
"01110110", 
"01010001", 
"10010000", 
"01110011", 
"01110111", 
"01100100", 
"01010110", 
"10000110", 
"01111101", 
"10110011", 
"10010001", 
"10011111", 
"01111100", 
"01101011", 
"10001010", 
"01101111", 
"01001111", 
"10000101", 
"10011001", 
"10001101", 
"10000000", 
"01100011", 
"00111110", 
"01111111", 
"01111000", 
"01011010", 
"01100100", 
"10101111", 
"10101001", 
"01100110", 
"10000111", 
"10000110", 
"01110010", 
"01011100", 
"10000110", 
"01110100", 
"10010001", 
"01001010", 
"10010101", 
"10000010", 
"01100111", 
"10110100", 
"01000111", 
"01110000", 
"10101110", 
"01011101", 
"01101111", 
"01111010", 
"01101001", 
"10000110", 
"01100011", 
"01101101", 
"01100111", 
"01011101", 
"01100111", 
"01000111", 
"10000011", 
"10100000", 
"01110110", 
"01010100", 
"10011111", 
"01011001", 
"01101000", 
"01111100", 
"01100111", 
"01101010", 
"10100001", 
"01100100", 
"01110101", 
"01111010", 
"01100001", 
"10000011", 
"01101000", 
"10001011", 
"10010000", 
"01010101", 
"10111101", 
"01110011", 
"10000110", 
"10001011", 
"01001100", 
"01101111", 
"01101110", 
"01100001", 
"10001011", 
"01101110", 
"01000001", 
"01100010", 
"01110111", 
"10011110", 
"01110011", 
"01111111", 
"10101001", 
"01101001", 
"01101001", 
"01110010", 
"10000101", 
"01111011", 
"10010001", 
"10101011", 
"01010110", 
"01101000", 
"01011100", 
"01111010", 
"01101001", 
"01110100", 
"10000011", 
"01010010", 
"10011011", 
"01100011", 
"10000011", 
"10001100", 
"01110100", 
"01101110", 
"01101101", 
"01011101", 
"01101110", 
"01110100", 
"01010011", 
"10100111", 
"01101101", 
"01110101", 
"01010011", 
"01110010", 
"10001001", 
"01011011", 
"10000100", 
"01101010", 
"01010110", 
"01011110", 
"00110100", 
"01011111", 
"01111010", 
"01101001", 
"01111100", 
"01111001", 
"01111110", 
"01011110", 
"10000100", 
"10101011", 
"01010001", 
"01110101", 
"01101100", 
"10001010", 
"01010100", 
"01101111", 
"10001010", 
"10011110", 
"10000001", 
"01000001", 
"01101101", 
"01010010", 
"01110101", 
"01010101", 
"01010000", 
"11001101", 
"01110001", 
"10000110", 
"10001100", 
"01111100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_51: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_51(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
