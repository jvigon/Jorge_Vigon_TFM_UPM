use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_39_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_39_LAYER;

architecture Behavioral of ROM_FC_120_39_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_39: ROM_ARRAY_PESOS_FC_120 := (
"10100100", 
"10011001", 
"10101100", 
"01111101", 
"01010100", 
"01000001", 
"10000100", 
"10001110", 
"01110010", 
"01110001", 
"10000000", 
"00011010", 
"01101111", 
"11001001", 
"10010110", 
"10100101", 
"01110010", 
"01101101", 
"01100011", 
"01001110", 
"01111001", 
"01001110", 
"01101001", 
"01101111", 
"11000101", 
"10100001", 
"01111000", 
"01110100", 
"01101000", 
"10101010", 
"01111001", 
"10011110", 
"10011100", 
"01111010", 
"10000100", 
"10001011", 
"10001111", 
"01111011", 
"01001101", 
"01111011", 
"10001110", 
"10001110", 
"00110100", 
"10010100", 
"10001001", 
"01110100", 
"01110101", 
"10001100", 
"01111101", 
"01110100", 
"10001001", 
"01110110", 
"10000100", 
"10011110", 
"01110010", 
"01100100", 
"10011011", 
"01001100", 
"00111110", 
"01101010", 
"10010000", 
"10000100", 
"10000101", 
"01110011", 
"10000010", 
"11000110", 
"01111010", 
"01100000", 
"10101101", 
"11000100", 
"10000010", 
"01110011", 
"01101011", 
"10000011", 
"10101111", 
"01100010", 
"10101011", 
"01010001", 
"01101111", 
"01111100", 
"10010110", 
"01110001", 
"01101100", 
"01000011", 
"10111101", 
"10011101", 
"01111111", 
"01100010", 
"10000100", 
"10010001", 
"10101000", 
"01101001", 
"01110100", 
"01011000", 
"01101111", 
"01110111", 
"01110100", 
"10010111", 
"10010010", 
"01011000", 
"01111000", 
"01111001", 
"10001010", 
"00111010", 
"01011100", 
"10101101", 
"01110011", 
"10011100", 
"01111110", 
"01111100", 
"01100011", 
"10000011", 
"10001011", 
"10101110", 
"01001010", 
"01110010", 
"10000110", 
"10001111", 
"01000010", 
"01001000", 
"10011001", 
"01111010", 
"01111111", 
"10001110", 
"10011011", 
"01111000", 
"10001111", 
"01111011", 
"10000101", 
"01111101", 
"01100101", 
"01011011", 
"10010001", 
"10100100", 
"01001100", 
"10100100", 
"01101100", 
"10010111", 
"10001001", 
"01110101", 
"01101010", 
"10011011", 
"01101011", 
"01111010", 
"01011010", 
"01011001", 
"00110111", 
"01110001", 
"10010000", 
"10100100", 
"10011010", 
"10011010", 
"01011000", 
"00110111", 
"01100001", 
"01111011", 
"01000011", 
"10101001", 
"01011100", 
"10001000", 
"10101111", 
"01111011", 
"01111011", 
"10010100", 
"10010000", 
"10001101", 
"11001110", 
"01010100", 
"10001001", 
"01100100", 
"01010100", 
"10101110", 
"01111100", 
"01101010", 
"10000011", 
"01100010", 
"10111010", 
"10001000", 
"01111110", 
"10000011", 
"10001100", 
"10010001", 
"10010011", 
"01010010", 
"10101101", 
"01010010", 
"10000111", 
"10011001", 
"01101111", 
"01011110", 
"01101111", 
"01110101", 
"01100110", 
"01110110", 
"00011111", 
"00111001", 
"10010101", 
"10000010", 
"01110110", 
"11100000", 
"10001011", 
"01011010", 
"01010000", 
"01001000", 
"01010100", 
"10011001", 
"01111000", 
"01101011", 
"10010000", 
"01011110", 
"01100011", 
"01011110", 
"10001110", 
"01101100", 
"01111011", 
"10000011", 
"01111000", 
"00100111", 
"00111010", 
"01111100", 
"00101011", 
"01101010", 
"10001011", 
"01100001", 
"10001100", 
"00101100", 
"10011001", 
"10001011", 
"10100011", 
"10101011", 
"10011101", 
"00101101", 
"10001010", 
"01111101", 
"01111101", 
"01110100", 
"01111111", 
"00001101", 
"01111000", 
"10000110", 
"10001111", 
"01111111", 
"01100101", 
"10110100", 
"10000001", 
"01010011", 
"01100001", 
"10010001", 
"10011011", 
"10010010", 
"10100001", 
"00110101", 
"01101000", 
"01101000", 
"10001011", 
"01110101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_39: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_39(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
