use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_71_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_71_LAYER;

architecture Behavioral of ROM_FC_120_71_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_71: ROM_ARRAY_PESOS_FC_120 := (
"01100100", 
"10100011", 
"10000010", 
"01111100", 
"01110001", 
"01111000", 
"10011000", 
"10010001", 
"01111000", 
"01010011", 
"10001111", 
"00100011", 
"01001010", 
"01010010", 
"10010101", 
"10001001", 
"01111001", 
"01110000", 
"10001001", 
"01111001", 
"01010001", 
"01110011", 
"10110110", 
"10111001", 
"10000100", 
"10000111", 
"10111011", 
"00000000", 
"10001011", 
"01010011", 
"10001110", 
"01111110", 
"10001100", 
"00101011", 
"01111101", 
"01111100", 
"01100100", 
"00101111", 
"10001000", 
"01111011", 
"01111000", 
"10101100", 
"01111010", 
"01001010", 
"10001100", 
"01101000", 
"01111011", 
"01110110", 
"01110110", 
"00010011", 
"10100010", 
"10011101", 
"01111000", 
"01010000", 
"01000101", 
"10011110", 
"01110111", 
"10111010", 
"10010111", 
"10001011", 
"10011000", 
"00111010", 
"10001011", 
"01101011", 
"10000001", 
"01000000", 
"10011001", 
"01111110", 
"01100111", 
"01001011", 
"01101001", 
"01010001", 
"10000010", 
"10110010", 
"01111001", 
"01001000", 
"01011110", 
"01110101", 
"10001010", 
"01101110", 
"10011111", 
"01101010", 
"01111001", 
"01110000", 
"10000011", 
"10100011", 
"01111001", 
"01011110", 
"10011001", 
"10010000", 
"10100001", 
"01101001", 
"01101011", 
"10000011", 
"10001000", 
"10000100", 
"10100011", 
"01111100", 
"01100111", 
"10000011", 
"01110100", 
"01100110", 
"10001000", 
"01111010", 
"10000110", 
"10000101", 
"10011111", 
"01101111", 
"01000111", 
"10110101", 
"10010100", 
"10010011", 
"01000001", 
"01011000", 
"01011100", 
"01000001", 
"01101110", 
"01100111", 
"01101010", 
"01010011", 
"01110110", 
"10100000", 
"10000101", 
"10110100", 
"10101000", 
"11000001", 
"10001000", 
"10010001", 
"01111011", 
"01101111", 
"10010101", 
"10000111", 
"01110011", 
"01111011", 
"00110001", 
"10100001", 
"01110111", 
"10100100", 
"01011111", 
"01110001", 
"10000011", 
"01110100", 
"10001011", 
"10000000", 
"10000100", 
"01001101", 
"10001101", 
"10001110", 
"01110001", 
"10011010", 
"01111011", 
"10110010", 
"10000101", 
"01110101", 
"10000010", 
"10001011", 
"10001000", 
"10100111", 
"01110100", 
"01111001", 
"01101010", 
"10110000", 
"10000010", 
"10001010", 
"01111100", 
"01010010", 
"10010001", 
"01101000", 
"01110010", 
"01011011", 
"01110000", 
"10001010", 
"01100000", 
"11001001", 
"10000100", 
"01101110", 
"10001101", 
"11000111", 
"10001101", 
"00110011", 
"01110000", 
"10100101", 
"10001110", 
"00111100", 
"01110010", 
"00111101", 
"01111101", 
"10111000", 
"11000101", 
"10100100", 
"01101001", 
"10011010", 
"10001001", 
"10011101", 
"10010000", 
"01100000", 
"10010001", 
"01010101", 
"01011100", 
"10110110", 
"10001010", 
"10000111", 
"01110101", 
"01111010", 
"10010101", 
"10001110", 
"01110111", 
"01111110", 
"10010010", 
"10101111", 
"10000010", 
"10010000", 
"01101101", 
"01100011", 
"01110110", 
"10011001", 
"10001001", 
"10000000", 
"10001110", 
"01101110", 
"10101111", 
"10001011", 
"01111111", 
"10000100", 
"10000000", 
"10101011", 
"10000101", 
"01100100", 
"10010001", 
"10010010", 
"10010011", 
"01110100", 
"01111110", 
"10011110", 
"01101100", 
"01111111", 
"10101110", 
"10101001", 
"10011001", 
"10010111", 
"10100110", 
"10110000", 
"10001110", 
"00100101", 
"10010000", 
"10001001", 
"01010000", 
"01111001", 
"01111111", 
"10011000", 
"01101011", 
"01110110", 
"10100100", 
"01110010", 
"10010001", 
"01101111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_71: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_71(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
