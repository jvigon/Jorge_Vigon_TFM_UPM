use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_82_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_82_LAYER;

architecture Behavioral of ROM_FC_84_82_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_82: ROM_ARRAY_PESOS_FC_84 := (
"10011011", 
"01101000", 
"01101110", 
"10011010", 
"10010010", 
"10000111", 
"01111011", 
"01001001", 
"01010110", 
"01111000", 
"10001100", 
"10101011", 
"10001101", 
"10010000", 
"10010110", 
"01111110", 
"10011001", 
"01101001", 
"10010011", 
"01000100", 
"10010100", 
"00100111", 
"01101100", 
"01100111", 
"01110110", 
"01101111", 
"01010000", 
"01101000", 
"10101001", 
"10011100", 
"01110100", 
"10000110", 
"01101101", 
"01100000", 
"01101100", 
"01101011", 
"01111000", 
"10100001", 
"01010111", 
"10011000", 
"10010100", 
"10000100", 
"10101111", 
"01001000", 
"10010010", 
"01111001", 
"10101011", 
"10011100", 
"10000100", 
"01111101", 
"10000111", 
"01111010", 
"01101011", 
"10001110", 
"01001100", 
"10010100", 
"10010011", 
"01111101", 
"10010100", 
"10000000", 
"10001100", 
"01001111", 
"01111101", 
"00111111", 
"10001111", 
"01101100", 
"10011001", 
"10000001", 
"10010101", 
"01100100", 
"10000100", 
"01111110", 
"01010100", 
"01100000", 
"10011010", 
"10000101", 
"01100000", 
"10000111", 
"10011110", 
"10000010", 
"01110001", 
"10000101", 
"01100110", 
"10011110", 
"10100001", 
"10010111", 
"10101101", 
"10011000", 
"01101011", 
"10110000", 
"01111111", 
"01100000", 
"10100000", 
"10010011", 
"01010001", 
"01110110", 
"10000001", 
"10010011", 
"01010110", 
"10001001", 
"01111101", 
"10101100", 
"10001011", 
"01011011", 
"10100101", 
"10011001", 
"01011111", 
"01101111", 
"10010010", 
"01001000", 
"10000010", 
"10000011", 
"01101101", 
"01001110", 
"01110110", 
"01111110", 
"01110101", 
"01000011", 
"10000110", 
"01001101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_82: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_82(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
