use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_73_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_73_LAYER;

architecture Behavioral of ROM_FC_120_73_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_73: ROM_ARRAY_PESOS_FC_120 := (
"10000001", 
"01111110", 
"10001111", 
"01101000", 
"01111100", 
"01001001", 
"01110111", 
"01101110", 
"01101010", 
"10001011", 
"01111001", 
"10001000", 
"10011001", 
"00111110", 
"10000010", 
"10010001", 
"01111000", 
"01100111", 
"01111101", 
"01010100", 
"10000011", 
"10001110", 
"01100101", 
"01011101", 
"01101111", 
"01111110", 
"10010001", 
"10101001", 
"10010001", 
"01011111", 
"01101000", 
"01111001", 
"10001100", 
"10010000", 
"10010111", 
"01001111", 
"01110011", 
"10000001", 
"00100110", 
"01101000", 
"10000010", 
"01110111", 
"01110101", 
"10010110", 
"01111011", 
"10111000", 
"01111110", 
"10001011", 
"01101111", 
"10010101", 
"01000110", 
"01101100", 
"10000111", 
"10000000", 
"01010001", 
"01101101", 
"01101110", 
"00100000", 
"01100111", 
"10010110", 
"01011100", 
"11000001", 
"01110110", 
"01110110", 
"10010000", 
"01110000", 
"01101001", 
"10001100", 
"01111100", 
"00001000", 
"10010110", 
"10100001", 
"10001110", 
"10000010", 
"10000010", 
"01110010", 
"10101000", 
"10000001", 
"10001000", 
"01111010", 
"10001101", 
"10000011", 
"10010001", 
"10001110", 
"10011101", 
"10001000", 
"01110100", 
"10000010", 
"01110111", 
"01010000", 
"01101100", 
"01111001", 
"01110011", 
"10001100", 
"01101001", 
"10010010", 
"10010011", 
"10000101", 
"10010000", 
"10100101", 
"01111011", 
"01111101", 
"01111000", 
"01110110", 
"01101011", 
"10000100", 
"01100101", 
"10011101", 
"10000001", 
"10011010", 
"01101011", 
"01101111", 
"10100001", 
"10100110", 
"01110110", 
"01000100", 
"01110001", 
"01101001", 
"10001000", 
"01100101", 
"10001000", 
"01100111", 
"01011100", 
"10010111", 
"10110001", 
"01111011", 
"01101111", 
"10001100", 
"01011100", 
"10110100", 
"10111010", 
"01010001", 
"10100010", 
"01000010", 
"10100101", 
"10000100", 
"10000010", 
"01111001", 
"01111110", 
"10001100", 
"10111100", 
"01011011", 
"01111010", 
"01101110", 
"01110100", 
"10100011", 
"01111010", 
"01101010", 
"10001010", 
"10010000", 
"01110000", 
"01101010", 
"01110110", 
"10010000", 
"01101001", 
"01110000", 
"10100001", 
"01000010", 
"01111100", 
"10000111", 
"10001000", 
"10011011", 
"01110101", 
"10001110", 
"10000110", 
"01010100", 
"01001111", 
"10101111", 
"01110010", 
"10100101", 
"01101110", 
"01110010", 
"10001000", 
"10001101", 
"01101010", 
"10000101", 
"10011001", 
"01100000", 
"01001000", 
"01111011", 
"10001111", 
"01011110", 
"01111011", 
"10010011", 
"10000101", 
"10010111", 
"01011000", 
"10000111", 
"10010111", 
"01000110", 
"10000011", 
"10001110", 
"01111000", 
"01110010", 
"01010001", 
"10010000", 
"01111110", 
"01000111", 
"01011110", 
"01111100", 
"01111100", 
"10100010", 
"10011011", 
"01110110", 
"01000111", 
"10100010", 
"10000010", 
"01111100", 
"00111101", 
"10001001", 
"10010000", 
"10000101", 
"01110110", 
"01100001", 
"10011010", 
"01111001", 
"10001110", 
"10001100", 
"01110111", 
"01010110", 
"01001111", 
"01111000", 
"01111101", 
"10001101", 
"01011100", 
"10010010", 
"10110011", 
"11001101", 
"01101111", 
"01110101", 
"01110010", 
"01000101", 
"10000010", 
"10000100", 
"01010100", 
"10101010", 
"01101011", 
"01011100", 
"10001100", 
"10001000", 
"01100110", 
"10000010", 
"10111111", 
"11011110", 
"10000011", 
"01001000", 
"01001111", 
"01010010", 
"10001100", 
"10101110", 
"00111011", 
"10111101", 
"10011001", 
"10100101", 
"01110110", 
"10000110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_73: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_73(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
