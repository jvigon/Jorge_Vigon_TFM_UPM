use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_29_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_29_LAYER;

architecture Behavioral of ROM_FC_120_29_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_29: ROM_ARRAY_PESOS_FC_120 := (
"10011011", 
"10100000", 
"10000110", 
"10101011", 
"01110011", 
"11011110", 
"01010100", 
"10000000", 
"01100100", 
"00110010", 
"01011100", 
"00111111", 
"01000010", 
"01110010", 
"01111111", 
"01101000", 
"10010110", 
"01110101", 
"01100000", 
"10110101", 
"10000110", 
"10110110", 
"10110011", 
"01110000", 
"10010011", 
"01000100", 
"01010111", 
"01010100", 
"01000000", 
"10100101", 
"10000111", 
"01110001", 
"10001110", 
"01001001", 
"01010111", 
"10100100", 
"10001000", 
"10010111", 
"10101000", 
"01110000", 
"10001000", 
"01100111", 
"10000100", 
"01100000", 
"01011001", 
"10000110", 
"01111011", 
"01111011", 
"10010111", 
"01011010", 
"10011101", 
"11000110", 
"10010001", 
"10011101", 
"10000000", 
"01111111", 
"01101001", 
"10000000", 
"10010011", 
"01101100", 
"01111111", 
"10010011", 
"10001000", 
"01101110", 
"01100101", 
"10010110", 
"10101101", 
"01110100", 
"10010110", 
"01101100", 
"01111001", 
"01110110", 
"10000011", 
"01110000", 
"10100001", 
"01000010", 
"01110101", 
"10110010", 
"10000101", 
"01111011", 
"01111000", 
"01111100", 
"10010001", 
"01011100", 
"10010001", 
"10000110", 
"10000110", 
"01011001", 
"10000010", 
"01111000", 
"01001111", 
"01011100", 
"10000000", 
"01110010", 
"10001010", 
"10000011", 
"10110110", 
"01110011", 
"10001111", 
"01111011", 
"01111100", 
"10010111", 
"01111100", 
"01011000", 
"10000110", 
"01110000", 
"10010011", 
"01011010", 
"01100110", 
"01011011", 
"10010010", 
"01110010", 
"10000011", 
"10000001", 
"10001101", 
"10000011", 
"01111010", 
"10011001", 
"10110111", 
"01110000", 
"01111101", 
"01110010", 
"10001110", 
"01110100", 
"01001100", 
"10011110", 
"10000101", 
"10000010", 
"01110010", 
"10011101", 
"01010001", 
"01111110", 
"10000101", 
"01011011", 
"10010110", 
"10010011", 
"10001111", 
"10101010", 
"10010000", 
"10001000", 
"01011011", 
"01100100", 
"01110111", 
"01100111", 
"10100111", 
"01011001", 
"01110001", 
"01000101", 
"10000110", 
"10110001", 
"01101000", 
"01011110", 
"10000110", 
"10110011", 
"10010011", 
"01101101", 
"01001101", 
"10111001", 
"01111011", 
"01111101", 
"10010001", 
"01100011", 
"01011000", 
"01011010", 
"10000100", 
"10010010", 
"01101011", 
"10100111", 
"10001011", 
"01111001", 
"10000000", 
"00111110", 
"01101110", 
"10011011", 
"01110000", 
"01110010", 
"01110000", 
"01000110", 
"01100001", 
"01110010", 
"10000110", 
"10101101", 
"01011000", 
"10001001", 
"01110001", 
"01011101", 
"10100001", 
"01111101", 
"01000110", 
"10001100", 
"10001100", 
"01111000", 
"10100100", 
"10000001", 
"01111100", 
"10010010", 
"10001111", 
"10101010", 
"01110111", 
"01101101", 
"01101000", 
"01101001", 
"01101100", 
"10000001", 
"10011110", 
"01011100", 
"10000101", 
"10000110", 
"10111010", 
"01011111", 
"01100101", 
"01100010", 
"01101101", 
"10110010", 
"00110101", 
"10001100", 
"10000011", 
"01011100", 
"10100111", 
"10010000", 
"10001011", 
"01011100", 
"01100111", 
"01111110", 
"01100010", 
"01101000", 
"01111110", 
"10100001", 
"10001001", 
"01011001", 
"01110110", 
"10010001", 
"01101100", 
"01001101", 
"10001010", 
"01101111", 
"10100111", 
"10010010", 
"01100010", 
"01111010", 
"01101110", 
"01101001", 
"01101000", 
"10101111", 
"01101011", 
"10010000", 
"01111101", 
"01000101", 
"01111101", 
"00110111", 
"01111100", 
"01011111", 
"01011100", 
"10101010", 
"01111110", 
"01110100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_29: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_29(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
