use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_70_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_70_LAYER;

architecture Behavioral of ROM_FC_84_70_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_70: ROM_ARRAY_PESOS_FC_84 := (
"01101110", 
"10010100", 
"01110111", 
"01101101", 
"01101000", 
"10001111", 
"01111111", 
"01111001", 
"01101011", 
"01111110", 
"01110001", 
"01010101", 
"10011101", 
"10011011", 
"01010110", 
"10011011", 
"10000010", 
"01110100", 
"10011010", 
"10000100", 
"01100000", 
"10000010", 
"10000000", 
"01100111", 
"10001101", 
"10001100", 
"10001001", 
"01100001", 
"01010101", 
"01111110", 
"10010001", 
"01011010", 
"10000000", 
"10000100", 
"01010000", 
"01110010", 
"01111010", 
"01100011", 
"01101110", 
"10001010", 
"10000000", 
"01110100", 
"01001101", 
"01110000", 
"01110011", 
"10010010", 
"01011000", 
"01111010", 
"01110001", 
"01100011", 
"01111111", 
"10001011", 
"10001000", 
"10010010", 
"10000110", 
"01010111", 
"01111001", 
"01101110", 
"01110110", 
"01100010", 
"01101010", 
"10001010", 
"10000100", 
"01110101", 
"10010111", 
"10101101", 
"10101111", 
"10001111", 
"10000100", 
"10011110", 
"01110010", 
"01101010", 
"10000100", 
"01011011", 
"01111101", 
"10000011", 
"01101011", 
"01110111", 
"01101111", 
"01101101", 
"10000111", 
"01100100", 
"10010001", 
"10011111", 
"01000001", 
"10001001", 
"10001011", 
"01001010", 
"01101000", 
"01100111", 
"01010000", 
"10001101", 
"10011011", 
"01101110", 
"01110111", 
"10010011", 
"10000001", 
"10001001", 
"10000100", 
"10100001", 
"10001100", 
"10010100", 
"01110000", 
"01110011", 
"01110011", 
"01100110", 
"01110001", 
"01110111", 
"01100110", 
"10001111", 
"01111110", 
"10010100", 
"01110011", 
"10000011", 
"10000010", 
"01110100", 
"01101110", 
"01011111", 
"01101001", 
"01010010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_70: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_70(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
