use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_55_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_55_LAYER;

architecture Behavioral of ROM_FC_84_55_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_55: ROM_ARRAY_PESOS_FC_84 := (
"01101101", 
"10000011", 
"01011111", 
"01100001", 
"10001011", 
"01100101", 
"01111001", 
"01001000", 
"10001100", 
"01101110", 
"10000100", 
"01101111", 
"01010111", 
"10110001", 
"01101100", 
"01010110", 
"01101010", 
"01101101", 
"10000010", 
"10000111", 
"10000110", 
"01011111", 
"01101110", 
"01111101", 
"10010001", 
"10111101", 
"01100011", 
"01111000", 
"01111001", 
"01010001", 
"01111110", 
"01111110", 
"01111110", 
"01111100", 
"01100111", 
"01100011", 
"01110010", 
"10000001", 
"10001010", 
"10000011", 
"01001101", 
"11001101", 
"01111011", 
"01110110", 
"01101110", 
"01000010", 
"01101001", 
"01100100", 
"01100010", 
"01111101", 
"10000101", 
"10010011", 
"10010110", 
"01001110", 
"10000000", 
"10011010", 
"10000001", 
"01110000", 
"01110111", 
"10001000", 
"01110010", 
"10001001", 
"01101101", 
"01111011", 
"10001100", 
"01101000", 
"01111011", 
"10001111", 
"01110101", 
"01100100", 
"01111100", 
"01111011", 
"01100111", 
"00111101", 
"01100110", 
"10000101", 
"01101000", 
"01101101", 
"01011010", 
"01100000", 
"01101110", 
"00111110", 
"01010001", 
"01100101", 
"01110110", 
"10001011", 
"01100101", 
"01100101", 
"01100001", 
"01011101", 
"10001001", 
"10011001", 
"01110101", 
"10000011", 
"01101000", 
"10011011", 
"01011110", 
"10000111", 
"10001100", 
"01110101", 
"01101111", 
"01100001", 
"01101001", 
"01111110", 
"01110001", 
"10010100", 
"10010110", 
"10000010", 
"10000100", 
"01111100", 
"10000010", 
"10011001", 
"10011000", 
"01101000", 
"01101110", 
"10001010", 
"01100011", 
"10100101", 
"10010100", 
"10000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_55: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_55(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
