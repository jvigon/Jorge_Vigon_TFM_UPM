use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_117_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_117_LAYER;

architecture Behavioral of ROM_FC_120_117_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_117: ROM_ARRAY_PESOS_FC_120 := (
"10101001", 
"01110001", 
"00111010", 
"10101110", 
"10000001", 
"11001001", 
"01111000", 
"01000010", 
"01011000", 
"10001110", 
"10010011", 
"01110111", 
"01001100", 
"01011011", 
"01110010", 
"10000010", 
"10101110", 
"00110000", 
"01101100", 
"11000100", 
"10010100", 
"10111010", 
"01101111", 
"11000011", 
"01110100", 
"01111000", 
"01111010", 
"01010110", 
"00100100", 
"01101011", 
"01101001", 
"10011001", 
"10111011", 
"01100111", 
"01110100", 
"01111000", 
"10100100", 
"01111000", 
"10110110", 
"11001010", 
"01010101", 
"00111111", 
"01110000", 
"10001001", 
"01101101", 
"01101001", 
"01110101", 
"10000100", 
"01111111", 
"01011000", 
"01110111", 
"00110000", 
"01110010", 
"00111100", 
"10000011", 
"10001001", 
"10000111", 
"00000110", 
"00111111", 
"10010011", 
"10111110", 
"01101001", 
"01100110", 
"10001011", 
"01110011", 
"01011011", 
"01101101", 
"01111001", 
"01010000", 
"10010000", 
"01110010", 
"01101000", 
"10010100", 
"01100101", 
"01100110", 
"01001111", 
"01000010", 
"10111100", 
"01111001", 
"01111010", 
"01001001", 
"00000000", 
"10100011", 
"01111111", 
"10000010", 
"10011001", 
"10111101", 
"01111011", 
"01010000", 
"01111101", 
"01111111", 
"01011001", 
"01000010", 
"10111010", 
"01111101", 
"01110011", 
"01110101", 
"01011001", 
"10011010", 
"10001011", 
"10101101", 
"01010111", 
"10011111", 
"10011100", 
"00111010", 
"11001011", 
"01110011", 
"01010000", 
"11100010", 
"10101011", 
"01101001", 
"10001001", 
"00011110", 
"10101100", 
"11100001", 
"00101011", 
"10101101", 
"01001110", 
"01100101", 
"01011101", 
"01101010", 
"10000111", 
"01101100", 
"01111110", 
"11010101", 
"10011001", 
"01110101", 
"10100001", 
"01100101", 
"10010011", 
"10010000", 
"10001010", 
"01011010", 
"10001110", 
"01111101", 
"01001001", 
"10001111", 
"01001110", 
"01101100", 
"01001100", 
"01110000", 
"11001000", 
"10000011", 
"10000001", 
"01100101", 
"01100010", 
"01111010", 
"01111010", 
"10000100", 
"01010110", 
"01100101", 
"01011101", 
"01111000", 
"01001110", 
"10011001", 
"01101111", 
"01011011", 
"01110010", 
"10000111", 
"10010101", 
"01010101", 
"01010000", 
"10001100", 
"10110101", 
"10000100", 
"01001010", 
"10000011", 
"01110001", 
"01110001", 
"10011111", 
"10011011", 
"01000110", 
"10000011", 
"01100001", 
"10001100", 
"10010000", 
"01011110", 
"10110011", 
"10110011", 
"01111001", 
"01111111", 
"01001000", 
"01000110", 
"01100010", 
"01111001", 
"01111101", 
"01101010", 
"10010110", 
"01111100", 
"01101110", 
"01110010", 
"10010001", 
"10000010", 
"10011111", 
"01101101", 
"01001110", 
"01110011", 
"01010001", 
"01001001", 
"00101110", 
"01101101", 
"10001111", 
"01101111", 
"01100110", 
"01111011", 
"10100011", 
"01100011", 
"01101011", 
"01011011", 
"10000010", 
"01110010", 
"01111101", 
"01110000", 
"10100100", 
"10000011", 
"01101101", 
"01101100", 
"10100010", 
"01101111", 
"00111101", 
"10100110", 
"01001111", 
"01101100", 
"10000111", 
"01100111", 
"01110110", 
"10000100", 
"10001001", 
"01111100", 
"01101001", 
"01011001", 
"10010011", 
"01111110", 
"10101101", 
"01011101", 
"01011001", 
"01000011", 
"01111010", 
"01110100", 
"01111101", 
"01111000", 
"01110100", 
"01110010", 
"01111101", 
"01111000", 
"01101101", 
"10001011", 
"10010011", 
"01101010", 
"10001101", 
"10000001", 
"01111010", 
"01100011", 
"01111010", 
"01111011", 
"10001000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_117 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_117(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
