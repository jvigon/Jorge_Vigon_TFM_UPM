use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_17_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_17_LAYER;

architecture Behavioral of ROM_FC_120_17_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_17: ROM_ARRAY_PESOS_FC_120 := (
"01110010", 
"10001011", 
"01100010", 
"10001100", 
"01101101", 
"01101111", 
"10010110", 
"01010010", 
"10000001", 
"01110110", 
"10000101", 
"01010001", 
"01011011", 
"01101100", 
"01110011", 
"01101111", 
"01110111", 
"01110100", 
"10000000", 
"10001010", 
"01110001", 
"10011010", 
"10001100", 
"01111100", 
"10000001", 
"01101001", 
"10010100", 
"01011011", 
"01101110", 
"10010011", 
"01110001", 
"10000001", 
"01110011", 
"01011111", 
"01111000", 
"10011011", 
"01101101", 
"01101001", 
"01100010", 
"01110101", 
"10000111", 
"01110010", 
"10010100", 
"10000101", 
"01101110", 
"01110100", 
"01110010", 
"01110010", 
"01101100", 
"01011001", 
"01110111", 
"10001000", 
"01111000", 
"01111000", 
"10001111", 
"01110001", 
"01111001", 
"01100010", 
"01010111", 
"01100011", 
"10001111", 
"01111100", 
"01111001", 
"10001111", 
"01101101", 
"01101011", 
"01111100", 
"01110111", 
"01101101", 
"01101111", 
"01101011", 
"01010010", 
"10000000", 
"10001011", 
"01111100", 
"01100010", 
"01111111", 
"01110001", 
"01111011", 
"10010000", 
"01010101", 
"01110110", 
"01101100", 
"10001010", 
"01111110", 
"10011010", 
"01110101", 
"10011001", 
"01111110", 
"01111111", 
"10000010", 
"01111000", 
"01100100", 
"10000110", 
"01101011", 
"01111000", 
"01111010", 
"01111110", 
"10001000", 
"01111011", 
"01111101", 
"01100101", 
"10001011", 
"01101110", 
"01111000", 
"10001111", 
"10000010", 
"10001010", 
"01111111", 
"01110010", 
"01110000", 
"10010011", 
"01110010", 
"01111100", 
"01111011", 
"01100101", 
"10000101", 
"01100100", 
"10000111", 
"01110101", 
"01111110", 
"01010011", 
"01111000", 
"01110100", 
"01101001", 
"01100010", 
"10001010", 
"01111011", 
"10000001", 
"10000001", 
"01101000", 
"01100101", 
"10000110", 
"01010011", 
"01110011", 
"01101010", 
"01111101", 
"01111010", 
"01011101", 
"10001111", 
"01101010", 
"01111111", 
"01110100", 
"01110011", 
"01011001", 
"01110100", 
"01110110", 
"10000001", 
"01110111", 
"10001000", 
"01011110", 
"01100111", 
"01111001", 
"01110010", 
"01101010", 
"01101100", 
"01101100", 
"10011100", 
"10001111", 
"01111100", 
"01010001", 
"10000001", 
"10100011", 
"10001110", 
"01111101", 
"01110001", 
"10010101", 
"10010000", 
"01111000", 
"01111000", 
"01110111", 
"01101101", 
"01101001", 
"10000001", 
"10000001", 
"10000111", 
"01101110", 
"10000100", 
"01110010", 
"01110001", 
"10000101", 
"01110000", 
"10010000", 
"01111111", 
"01110010", 
"10011010", 
"01011111", 
"01100010", 
"01110111", 
"01110111", 
"10000010", 
"01111011", 
"01111111", 
"01111001", 
"10000001", 
"01111010", 
"10000100", 
"01100101", 
"01110101", 
"01100111", 
"10010011", 
"01101000", 
"01100000", 
"10001000", 
"01111101", 
"10011100", 
"01101110", 
"10000111", 
"01101011", 
"01100111", 
"01100011", 
"01110001", 
"10010000", 
"10001000", 
"01110000", 
"01111010", 
"01111110", 
"01100100", 
"01110000", 
"10000001", 
"01111110", 
"01111100", 
"01111110", 
"01110101", 
"10000111", 
"01101011", 
"01010101", 
"10010000", 
"10001011", 
"01110001", 
"01110101", 
"01110010", 
"01111101", 
"01100011", 
"01110000", 
"10010101", 
"01110111", 
"10000010", 
"01111111", 
"01110101", 
"01110101", 
"01111110", 
"10011111", 
"01111000", 
"01111100", 
"10000011", 
"01111001", 
"01100000", 
"01101001", 
"01101100", 
"01111110", 
"01111011", 
"10001011", 
"10000111", 
"01111110", 
"10000111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_17: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_17(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
