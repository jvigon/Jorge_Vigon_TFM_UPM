use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_30_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_30_LAYER;

architecture Behavioral of ROM_FC_84_30_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_30: ROM_ARRAY_PESOS_FC_84 := (
"01101111", 
"10001100", 
"01110110", 
"10010011", 
"01110010", 
"01111000", 
"01111110", 
"01110101", 
"01110010", 
"10010111", 
"10000100", 
"01100001", 
"01111010", 
"01101011", 
"10000110", 
"01110010", 
"01111100", 
"01110110", 
"01011000", 
"01101101", 
"10100011", 
"01111001", 
"10100000", 
"10000001", 
"10010000", 
"10001101", 
"01100011", 
"01011100", 
"01011100", 
"10001010", 
"10000101", 
"01001111", 
"01100111", 
"01110001", 
"01111001", 
"10000111", 
"01101110", 
"01111010", 
"01111010", 
"01100001", 
"01001010", 
"01110101", 
"01101000", 
"10000000", 
"01110001", 
"01001111", 
"01101010", 
"10010001", 
"10001111", 
"01100111", 
"01111110", 
"01110101", 
"10001001", 
"10000001", 
"01101110", 
"10001011", 
"10011000", 
"01110111", 
"01100011", 
"10010110", 
"01110111", 
"01111111", 
"01110001", 
"01011100", 
"01101100", 
"10000011", 
"01111011", 
"01110101", 
"10011111", 
"01001101", 
"10000110", 
"01100100", 
"01010110", 
"01110110", 
"10000011", 
"10011011", 
"01101001", 
"10010011", 
"01101100", 
"01111110", 
"01111111", 
"01011010", 
"01010111", 
"01111110", 
"01101010", 
"10000011", 
"01101011", 
"01100101", 
"10010000", 
"01110010", 
"01100000", 
"10001000", 
"10100001", 
"01111110", 
"10001011", 
"01100100", 
"10000101", 
"10011110", 
"01100101", 
"01101101", 
"10011100", 
"10001001", 
"01111001", 
"01100000", 
"01101001", 
"10001001", 
"01011110", 
"01101010", 
"01101100", 
"10100001", 
"10000010", 
"10001101", 
"01110001", 
"10000101", 
"10000010", 
"01111011", 
"01110100", 
"10101101", 
"10000000", 
"01110000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_30 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_30(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
