use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_59_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_59_LAYER;

architecture Behavioral of ROM_FC_120_59_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_59: ROM_ARRAY_PESOS_FC_120 := (
"01111010", 
"01110010", 
"01001101", 
"10000110", 
"01101111", 
"10011010", 
"01100001", 
"01001011", 
"01111000", 
"01000000", 
"01101110", 
"11000110", 
"01010111", 
"01110001", 
"01101110", 
"10100101", 
"10000001", 
"01110010", 
"01001100", 
"01110100", 
"01111001", 
"10010101", 
"01100111", 
"01100000", 
"10001010", 
"01100100", 
"01111110", 
"10111001", 
"01011101", 
"10000011", 
"10000100", 
"10001001", 
"01111111", 
"10000001", 
"01111001", 
"10011000", 
"01110100", 
"10011100", 
"10100010", 
"01011011", 
"10001111", 
"01101001", 
"10001011", 
"10001011", 
"01000111", 
"10101001", 
"10000011", 
"01100100", 
"01100110", 
"01100000", 
"01101000", 
"10101100", 
"01110011", 
"10010000", 
"10010001", 
"01011011", 
"10000101", 
"01011100", 
"01010101", 
"10000110", 
"01101111", 
"01101000", 
"01101110", 
"10000111", 
"01110101", 
"01101111", 
"00111110", 
"01111011", 
"10000011", 
"10100011", 
"01001111", 
"01111100", 
"01110000", 
"01110000", 
"01110111", 
"01111011", 
"01001011", 
"00110110", 
"01111010", 
"01110010", 
"01110110", 
"01100010", 
"01100100", 
"01001110", 
"01101000", 
"10001000", 
"10011000", 
"01101000", 
"01110000", 
"01000100", 
"01011000", 
"01101101", 
"01010001", 
"10001011", 
"01101011", 
"10000110", 
"01110111", 
"01100011", 
"01001100", 
"10010010", 
"01110100", 
"10000010", 
"01101110", 
"01010010", 
"01110011", 
"01010011", 
"01110001", 
"10000110", 
"10000101", 
"10111000", 
"01110000", 
"10000000", 
"01111010", 
"01001000", 
"01100111", 
"01000010", 
"10000010", 
"01010001", 
"10110000", 
"01010111", 
"10001001", 
"10100001", 
"01000010", 
"10000011", 
"01000101", 
"01110001", 
"10001000", 
"01101100", 
"10001000", 
"01111110", 
"01001100", 
"01100110", 
"01110000", 
"10011000", 
"10101011", 
"01111000", 
"10001000", 
"01100100", 
"01001111", 
"10000010", 
"10010001", 
"00111001", 
"10010000", 
"01101001", 
"10000000", 
"01001100", 
"01010110", 
"01010010", 
"10001111", 
"10000101", 
"10101001", 
"01100001", 
"01111010", 
"01101010", 
"10000010", 
"01011110", 
"01111001", 
"01111110", 
"01110001", 
"01110111", 
"01110001", 
"01010001", 
"01110100", 
"10001101", 
"01101110", 
"10100100", 
"10001010", 
"00111111", 
"10010001", 
"01100110", 
"10000001", 
"01111100", 
"01110001", 
"10000100", 
"10001100", 
"01110011", 
"01011001", 
"10000010", 
"10001011", 
"10000001", 
"01110011", 
"01010111", 
"11001010", 
"01000011", 
"01111110", 
"10010111", 
"01000111", 
"01111110", 
"01100100", 
"01101110", 
"01110101", 
"01100000", 
"10000011", 
"10000110", 
"10001100", 
"01101101", 
"10010010", 
"01110111", 
"10001110", 
"01100001", 
"10000001", 
"10010010", 
"10000100", 
"10010010", 
"10000101", 
"01010010", 
"01110101", 
"01101001", 
"01111000", 
"01110000", 
"10001100", 
"01101000", 
"01111100", 
"01111000", 
"01011001", 
"01110010", 
"10000001", 
"10011100", 
"01011011", 
"01001011", 
"01011100", 
"01100000", 
"01110110", 
"01111000", 
"10000011", 
"01111111", 
"01001000", 
"01101010", 
"10001000", 
"10000110", 
"10001001", 
"01110110", 
"10000010", 
"01101101", 
"10010001", 
"01011000", 
"01011100", 
"10101100", 
"01110010", 
"01110100", 
"01101100", 
"01001011", 
"10001000", 
"10001100", 
"01111011", 
"01010001", 
"11011010", 
"01011110", 
"01101001", 
"01000011", 
"01011101", 
"01110110", 
"10001101", 
"01101000", 
"01110111", 
"10000001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_59: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_59(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
