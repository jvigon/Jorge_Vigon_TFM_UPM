use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_63_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_63_LAYER;

architecture Behavioral of ROM_FC_120_63_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_63: ROM_ARRAY_PESOS_FC_120 := (
"10100100", 
"01111011", 
"00111111", 
"10100111", 
"10000011", 
"01100100", 
"01010111", 
"10000000", 
"10000101", 
"01000110", 
"00111110", 
"00111111", 
"00010101", 
"01110010", 
"01110100", 
"01110110", 
"10000111", 
"01100100", 
"01101110", 
"01001110", 
"10001001", 
"10000000", 
"10001101", 
"01111111", 
"01100101", 
"01010010", 
"01001101", 
"10010111", 
"01100110", 
"10110101", 
"01100010", 
"01100110", 
"01110101", 
"01010101", 
"10100110", 
"10010000", 
"01110110", 
"00110000", 
"01011011", 
"01011011", 
"01101000", 
"10011011", 
"10000100", 
"10000001", 
"10011101", 
"01000111", 
"01101011", 
"01100100", 
"01010001", 
"01111100", 
"11000011", 
"01100001", 
"01101100", 
"01001101", 
"01011001", 
"10000100", 
"01000111", 
"10111010", 
"01111011", 
"01111001", 
"10101010", 
"00010101", 
"10010100", 
"01110010", 
"10110001", 
"01111010", 
"01111101", 
"01011101", 
"01011111", 
"00111100", 
"01010011", 
"01101000", 
"10000111", 
"01100100", 
"00101001", 
"01110110", 
"01011111", 
"11001000", 
"01110001", 
"10000110", 
"01100001", 
"01111110", 
"10000101", 
"10001001", 
"01100110", 
"10000101", 
"10010010", 
"00001100", 
"01100110", 
"10000111", 
"01100010", 
"10010000", 
"10011101", 
"10010010", 
"10001001", 
"10001100", 
"00111101", 
"01101110", 
"01111110", 
"01101000", 
"01010010", 
"10010100", 
"01001011", 
"01000011", 
"01111001", 
"10101010", 
"10001100", 
"01100011", 
"10001110", 
"01101011", 
"01101011", 
"01110000", 
"01101101", 
"01111001", 
"10001011", 
"01110110", 
"01111100", 
"10000010", 
"01010001", 
"10011110", 
"01011011", 
"11010010", 
"01101011", 
"10010111", 
"01111010", 
"10000011", 
"01100110", 
"01111111", 
"10011010", 
"10101111", 
"10110101", 
"10010101", 
"01000101", 
"01111011", 
"01100100", 
"01101101", 
"10000100", 
"10011110", 
"01111110", 
"01100110", 
"10110101", 
"11010011", 
"01111011", 
"10001000", 
"01101101", 
"10000001", 
"10000111", 
"10001111", 
"10000100", 
"10011100", 
"01111111", 
"01101001", 
"10000000", 
"10010000", 
"01001111", 
"01011101", 
"10001011", 
"10101001", 
"01100011", 
"10010111", 
"10001101", 
"10010000", 
"01010110", 
"01110101", 
"01110101", 
"10001100", 
"10010000", 
"00111111", 
"01100001", 
"00111100", 
"10010101", 
"01011100", 
"01101001", 
"11001001", 
"10100011", 
"01111000", 
"10100011", 
"10001011", 
"01010000", 
"01010101", 
"01110111", 
"01110011", 
"01100110", 
"01101100", 
"00111010", 
"01000000", 
"10010001", 
"10010101", 
"01110110", 
"10100111", 
"10000001", 
"01110100", 
"01100100", 
"10110000", 
"10010100", 
"01011110", 
"10101010", 
"01001100", 
"01101110", 
"01010000", 
"01111011", 
"10010100", 
"10010001", 
"01110000", 
"10110110", 
"01101000", 
"01100010", 
"01111010", 
"01111111", 
"10100000", 
"10000111", 
"01110100", 
"10011101", 
"10010000", 
"01110000", 
"01111100", 
"01100011", 
"10100000", 
"01110011", 
"01010101", 
"10001101", 
"01110000", 
"10000000", 
"10000111", 
"10110110", 
"10001010", 
"01100110", 
"01111011", 
"10010010", 
"10000100", 
"10111001", 
"10010100", 
"01001010", 
"10001000", 
"01110011", 
"01010001", 
"00110101", 
"10111001", 
"01110011", 
"10010100", 
"10100111", 
"01101001", 
"01011101", 
"01101111", 
"10001111", 
"10000001", 
"10000001", 
"10010010", 
"01110111", 
"01011001", 
"01101100", 
"10001110", 
"01101010", 
"01110100", 
"10000000", 
"10010010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_63: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_63(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
