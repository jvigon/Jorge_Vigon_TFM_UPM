use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_28_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_28_LAYER;

architecture Behavioral of ROM_FC_120_28_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_28: ROM_ARRAY_PESOS_FC_120 := (
"10111000", 
"01101110", 
"01111100", 
"01010111", 
"10000010", 
"00100101", 
"01010101", 
"10001100", 
"01111100", 
"01101111", 
"01000011", 
"10001010", 
"01110001", 
"01011111", 
"10001000", 
"01111000", 
"01101100", 
"01100000", 
"10011101", 
"00111111", 
"10010101", 
"01010101", 
"01101000", 
"01010110", 
"10000010", 
"10010110", 
"01010111", 
"01111010", 
"01110101", 
"10001010", 
"10000110", 
"10000011", 
"01010110", 
"10001001", 
"10001111", 
"01101010", 
"10100000", 
"10100000", 
"01011100", 
"00111101", 
"01110000", 
"01110111", 
"01101110", 
"10001101", 
"01111100", 
"11000111", 
"10000001", 
"01110011", 
"01010110", 
"10001001", 
"01111100", 
"10100000", 
"01100101", 
"10001101", 
"01111000", 
"00101000", 
"10010001", 
"00010110", 
"01100111", 
"01100101", 
"01110010", 
"10111111", 
"10001111", 
"10001011", 
"10100011", 
"10011111", 
"10101110", 
"01011100", 
"01001011", 
"01001000", 
"10011110", 
"01111001", 
"01111011", 
"01110010", 
"10000000", 
"01111000", 
"11100010", 
"01111100", 
"10001011", 
"01110011", 
"01101101", 
"10011100", 
"01111110", 
"01101100", 
"10101110", 
"01011110", 
"01100110", 
"01110101", 
"01111110", 
"01101011", 
"01101100", 
"01101010", 
"10011010", 
"01100011", 
"10010101", 
"10000010", 
"01111100", 
"01110111", 
"10100110", 
"10000010", 
"01011010", 
"10001100", 
"01101101", 
"10001011", 
"01111100", 
"10000001", 
"01010011", 
"10000010", 
"01101101", 
"01111100", 
"10011001", 
"01111000", 
"01111010", 
"10000100", 
"10011100", 
"10000101", 
"01101000", 
"01010011", 
"10101010", 
"00111011", 
"01111111", 
"01101010", 
"01001111", 
"10100011", 
"10010111", 
"01011010", 
"10001010", 
"10000100", 
"10000010", 
"01110101", 
"10110011", 
"10010110", 
"10011010", 
"10000100", 
"10010001", 
"10001100", 
"10000101", 
"10001100", 
"10001000", 
"01010100", 
"10000001", 
"01110110", 
"10001000", 
"01101000", 
"01111101", 
"10000011", 
"10001000", 
"01011111", 
"10001100", 
"10011011", 
"01011000", 
"01111101", 
"10001100", 
"10010011", 
"01111100", 
"01101011", 
"10000110", 
"01111110", 
"01110011", 
"10001001", 
"10000100", 
"01100111", 
"10000000", 
"01111100", 
"10000111", 
"01011111", 
"01010111", 
"10010011", 
"01101101", 
"10010110", 
"01101110", 
"01110110", 
"10011001", 
"10010011", 
"01101101", 
"01110111", 
"10100000", 
"01110010", 
"10000000", 
"01101111", 
"01111110", 
"01001111", 
"01101101", 
"10010111", 
"10000011", 
"10111011", 
"01000111", 
"10100100", 
"10000010", 
"01100000", 
"01110110", 
"10011000", 
"10000111", 
"01100110", 
"10001011", 
"10110101", 
"01111110", 
"10000010", 
"01010010", 
"01110011", 
"10000011", 
"10100001", 
"10001100", 
"01001011", 
"00110001", 
"01100101", 
"01110000", 
"01111010", 
"01100000", 
"01110011", 
"10001001", 
"10011100", 
"01110011", 
"10010101", 
"10001110", 
"01111101", 
"10001110", 
"10001100", 
"10000000", 
"10000000", 
"01110101", 
"10010011", 
"01110100", 
"10000100", 
"01100101", 
"10000110", 
"10100100", 
"01011100", 
"01110100", 
"01011110", 
"01110001", 
"01101111", 
"10010011", 
"10101000", 
"01000101", 
"10011001", 
"10100011", 
"01110010", 
"01111100", 
"10000000", 
"01100100", 
"10011000", 
"01100100", 
"01011101", 
"01111001", 
"01001001", 
"01101010", 
"11001101", 
"01111110", 
"10110001", 
"00100100", 
"11000000", 
"01111100", 
"10001110", 
"10011100", 
"01111001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_28: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_28(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
