use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_55_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_55_LAYER;

architecture Behavioral of ROM_FC_120_55_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_55: ROM_ARRAY_PESOS_FC_120 := (
"10000111", 
"10000011", 
"10001000", 
"01001000", 
"01100101", 
"01011010", 
"10001011", 
"01101101", 
"10000110", 
"10010011", 
"10010111", 
"10010011", 
"01111000", 
"01010101", 
"01111110", 
"10000000", 
"01101101", 
"10000101", 
"10000110", 
"00101010", 
"01110001", 
"01001110", 
"01011100", 
"01110110", 
"01111011", 
"01101010", 
"01000111", 
"10001110", 
"01101101", 
"01101011", 
"10001101", 
"01111110", 
"01110100", 
"01101100", 
"01111101", 
"10110101", 
"01111011", 
"01110100", 
"01110100", 
"01100110", 
"10000010", 
"01111100", 
"01101011", 
"00111101", 
"01001010", 
"10011000", 
"01101100", 
"10001101", 
"01110100", 
"01011111", 
"01110000", 
"11010011", 
"10000011", 
"01001100", 
"10100010", 
"01101100", 
"10000101", 
"01010110", 
"01111101", 
"01111100", 
"01110000", 
"10011110", 
"10001010", 
"10000001", 
"01111001", 
"01101110", 
"01011010", 
"01101100", 
"01111011", 
"10000110", 
"01110111", 
"01001100", 
"01110011", 
"01101000", 
"01110101", 
"10100000", 
"10010001", 
"01100001", 
"10001010", 
"01110001", 
"10000010", 
"10000001", 
"01001101", 
"01011000", 
"10001000", 
"10010000", 
"01110001", 
"01011010", 
"10000001", 
"01101011", 
"01101110", 
"01110111", 
"01101101", 
"01110100", 
"10001001", 
"01110101", 
"01100101", 
"01001101", 
"01110010", 
"00111001", 
"10001000", 
"01101101", 
"01110010", 
"10000101", 
"10001001", 
"01110111", 
"01101110", 
"01101111", 
"01001111", 
"01111011", 
"01101110", 
"01101111", 
"01001100", 
"01110001", 
"01010001", 
"10001110", 
"01110001", 
"01100011", 
"10001101", 
"01100011", 
"01111111", 
"10000010", 
"01010110", 
"10000111", 
"01011011", 
"01011101", 
"10001010", 
"10000100", 
"01111110", 
"10000110", 
"10001001", 
"01110100", 
"10000110", 
"10101100", 
"01111100", 
"10000110", 
"10010001", 
"01100000", 
"01101000", 
"01101101", 
"00111010", 
"01110011", 
"10001100", 
"01110001", 
"01101101", 
"01010101", 
"01101000", 
"01101111", 
"10001010", 
"11001010", 
"10010001", 
"01110110", 
"01110100", 
"01110101", 
"01100110", 
"01110100", 
"01100010", 
"01110100", 
"10001000", 
"01111101", 
"01101001", 
"01100001", 
"01111010", 
"01100100", 
"01101110", 
"01000111", 
"01111000", 
"10010001", 
"01111101", 
"10010000", 
"01101110", 
"10101101", 
"10001010", 
"01011010", 
"10000101", 
"01111000", 
"10000001", 
"01100001", 
"01011110", 
"01000010", 
"01101001", 
"01101001", 
"10000011", 
"01110010", 
"10000101", 
"01111000", 
"01011111", 
"10100011", 
"10000000", 
"01010110", 
"10000100", 
"10001010", 
"01110000", 
"01110001", 
"01111010", 
"10010111", 
"10001010", 
"01101110", 
"01100100", 
"01010001", 
"10010001", 
"01100000", 
"01110000", 
"01100111", 
"01111101", 
"01010111", 
"01101110", 
"10001111", 
"10001000", 
"01110001", 
"01001000", 
"10000000", 
"01101101", 
"10011100", 
"01100100", 
"01010001", 
"01111101", 
"00111110", 
"10001101", 
"00100111", 
"10101011", 
"10000001", 
"01111111", 
"01111010", 
"01100100", 
"00110010", 
"01100110", 
"01111001", 
"10000110", 
"01011000", 
"01001000", 
"10000010", 
"01110011", 
"01011111", 
"01011001", 
"10000001", 
"10000101", 
"01101101", 
"01110100", 
"10001011", 
"01100100", 
"01010110", 
"01110100", 
"11000000", 
"10000000", 
"01000001", 
"01111101", 
"01000010", 
"01111010", 
"01110011", 
"01101010", 
"10001010", 
"10000011", 
"01100111", 
"01111101", 
"10001001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_55: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_55(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
