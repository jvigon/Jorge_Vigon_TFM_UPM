use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_66_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_66_LAYER;

architecture Behavioral of ROM_FC_120_66_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_66: ROM_ARRAY_PESOS_FC_120 := (
"10000000", 
"01001101", 
"01000111", 
"01011001", 
"01100110", 
"01101010", 
"01100011", 
"01101010", 
"10000100", 
"10011001", 
"01100010", 
"10001010", 
"01001111", 
"10100111", 
"10001101", 
"10000100", 
"01111010", 
"00010000", 
"01011001", 
"00111101", 
"01101000", 
"01101101", 
"01110111", 
"01101000", 
"01101001", 
"01110001", 
"01000101", 
"10110000", 
"01110010", 
"01001111", 
"10001010", 
"01111001", 
"01101111", 
"01011100", 
"01010001", 
"01001110", 
"10001001", 
"01110010", 
"01110001", 
"01001110", 
"01110101", 
"01100011", 
"01011011", 
"10011000", 
"10011110", 
"01111000", 
"01111001", 
"10000101", 
"01110101", 
"10010101", 
"01101111", 
"01010010", 
"10001000", 
"01100010", 
"01000101", 
"01110010", 
"10001101", 
"01101100", 
"01010101", 
"01111110", 
"10001000", 
"01101110", 
"10000101", 
"10010000", 
"01110100", 
"10000111", 
"01101011", 
"10000010", 
"10000101", 
"01100010", 
"10010010", 
"01110011", 
"01101010", 
"01101101", 
"01101101", 
"10001010", 
"10011011", 
"10001011", 
"10001100", 
"01101101", 
"01101110", 
"10000000", 
"01101010", 
"01101000", 
"01100011", 
"01010111", 
"01100000", 
"01110011", 
"01111101", 
"01111011", 
"01010110", 
"01101000", 
"01111011", 
"01110001", 
"01110111", 
"10001001", 
"01111011", 
"01101010", 
"01011000", 
"01101100", 
"01111010", 
"10000100", 
"01100001", 
"10010010", 
"01101010", 
"10101001", 
"01100001", 
"10001111", 
"10010010", 
"10000110", 
"01110110", 
"10000010", 
"10000110", 
"10000110", 
"01001101", 
"01111011", 
"01111111", 
"01011111", 
"10001101", 
"01101111", 
"10001101", 
"01100011", 
"01100001", 
"10101011", 
"01011010", 
"01001100", 
"10001100", 
"01111101", 
"10001011", 
"01100110", 
"01110010", 
"10000101", 
"10011000", 
"01111101", 
"10011001", 
"01011011", 
"10001000", 
"01001100", 
"01100011", 
"01100000", 
"10001010", 
"01110010", 
"01101110", 
"10001001", 
"01111000", 
"10011011", 
"01111111", 
"10011000", 
"10000010", 
"01111011", 
"00111110", 
"10100000", 
"10000111", 
"01111111", 
"01110001", 
"01100000", 
"01100010", 
"01111000", 
"01110110", 
"10000100", 
"01100011", 
"01110010", 
"01010111", 
"00110111", 
"10000100", 
"01011111", 
"00111000", 
"10100010", 
"01110011", 
"01110111", 
"01010010", 
"01110000", 
"01111001", 
"01110010", 
"01111010", 
"01110101", 
"01100101", 
"01001101", 
"01111101", 
"01110011", 
"01111000", 
"01010110", 
"01101111", 
"01111011", 
"10001001", 
"01101001", 
"01101000", 
"01111110", 
"01111001", 
"01111010", 
"01111101", 
"01101001", 
"01110110", 
"01100110", 
"10000100", 
"10011011", 
"10001110", 
"10000011", 
"01110110", 
"01100011", 
"01110101", 
"10010010", 
"01100011", 
"10000110", 
"01001100", 
"10001101", 
"10000000", 
"10000011", 
"01010000", 
"01101010", 
"01100100", 
"10000111", 
"10001110", 
"01000110", 
"10010000", 
"01110101", 
"10000110", 
"10011110", 
"01100110", 
"01110000", 
"01011011", 
"01010111", 
"01110101", 
"01101001", 
"01111000", 
"01001001", 
"01101101", 
"10001000", 
"01101001", 
"01000001", 
"00110111", 
"01101110", 
"01110011", 
"10001001", 
"01110101", 
"01101001", 
"01101000", 
"10000100", 
"01110111", 
"10000100", 
"01000111", 
"01001101", 
"01101100", 
"10001011", 
"10001000", 
"01100100", 
"01010111", 
"01100100", 
"10000010", 
"10010000", 
"01011011", 
"10010110", 
"10011110", 
"10001111", 
"01110110", 
"01101101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_66: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_66(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
