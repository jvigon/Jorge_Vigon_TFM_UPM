use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_75_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_75_LAYER;

architecture Behavioral of ROM_FC_84_75_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_75: ROM_ARRAY_PESOS_FC_84 := (
"10000000", 
"01011111", 
"01000000", 
"01110111", 
"10100110", 
"01101110", 
"10000011", 
"01101101", 
"10001000", 
"10001101", 
"01111001", 
"10001110", 
"10001001", 
"10100010", 
"01101101", 
"01110000", 
"10000001", 
"01110011", 
"01110100", 
"10010111", 
"00101100", 
"01101100", 
"01110100", 
"10001000", 
"10001001", 
"01110001", 
"10011000", 
"10011101", 
"10001011", 
"01011000", 
"01110010", 
"01110010", 
"01110001", 
"01101000", 
"01111100", 
"01000001", 
"10110011", 
"10000110", 
"10010111", 
"10010010", 
"01011111", 
"10011101", 
"10010110", 
"10000001", 
"01010000", 
"10001100", 
"01011111", 
"01101010", 
"10100001", 
"01110111", 
"10001101", 
"10011111", 
"01100101", 
"01111100", 
"10010100", 
"10111110", 
"10100001", 
"01111111", 
"01011111", 
"01111011", 
"10011001", 
"01000100", 
"01100111", 
"10110001", 
"01010101", 
"10000111", 
"01111101", 
"01100000", 
"10001001", 
"01111100", 
"01100101", 
"01111011", 
"01001101", 
"01111111", 
"10001000", 
"01111001", 
"10111011", 
"10001100", 
"01010011", 
"01010111", 
"10101110", 
"01011100", 
"01110111", 
"01111100", 
"10000100", 
"01011101", 
"01100011", 
"10010101", 
"10001101", 
"01111111", 
"01111011", 
"10011001", 
"10010100", 
"01010011", 
"10001110", 
"10110110", 
"10001000", 
"10010110", 
"01111001", 
"01100001", 
"10001001", 
"01101111", 
"01111111", 
"10000100", 
"10011001", 
"01111000", 
"10000111", 
"01110110", 
"01110101", 
"10001110", 
"00010011", 
"01111110", 
"01110100", 
"01011000", 
"01110101", 
"01010011", 
"01110111", 
"01100010", 
"10011101", 
"10101001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_75: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_75(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
