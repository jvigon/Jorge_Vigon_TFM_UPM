use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_65_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_65_LAYER;

architecture Behavioral of ROM_FC_84_65_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_65: ROM_ARRAY_PESOS_FC_84 := (
"01100101", 
"01111111", 
"01101001", 
"01101111", 
"10000001", 
"01110101", 
"10000101", 
"01011000", 
"01011011", 
"01101011", 
"10010001", 
"01111001", 
"01001110", 
"01111101", 
"01100100", 
"10010010", 
"10001000", 
"01011110", 
"10010001", 
"10001110", 
"10010001", 
"01100101", 
"01110001", 
"01111101", 
"01111011", 
"10010101", 
"01001001", 
"01101000", 
"10010000", 
"10010011", 
"10000000", 
"10000100", 
"01001000", 
"01101100", 
"01011110", 
"10000101", 
"01010110", 
"01101110", 
"01010100", 
"01011011", 
"01011100", 
"10010101", 
"01111101", 
"01010100", 
"01010101", 
"01010110", 
"10000010", 
"10010000", 
"10010000", 
"01101011", 
"01111010", 
"10101000", 
"01110110", 
"10001100", 
"01101100", 
"10100011", 
"10000111", 
"10001001", 
"10001010", 
"01111101", 
"10011010", 
"01110110", 
"01100011", 
"01000110", 
"11000100", 
"01010000", 
"10001111", 
"01100111", 
"10010110", 
"01011000", 
"10011100", 
"01110101", 
"01110001", 
"01110011", 
"01110111", 
"01101110", 
"10000100", 
"01110111", 
"10001010", 
"10010001", 
"01011101", 
"10000110", 
"01010000", 
"01111111", 
"01101101", 
"10000110", 
"10010101", 
"10001000", 
"01111001", 
"10110101", 
"01001001", 
"10000011", 
"01100000", 
"10111001", 
"01011100", 
"10001000", 
"10001001", 
"10000101", 
"10000000", 
"01110111", 
"01100101", 
"10000101", 
"10000000", 
"01010111", 
"10100111", 
"10010011", 
"10000101", 
"10001101", 
"01111110", 
"01110001", 
"01111101", 
"10100100", 
"10000011", 
"11000000", 
"01111011", 
"01111110", 
"01010100", 
"10110101", 
"01111101", 
"01100011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_65 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_65(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
