use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_81_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_81_LAYER;

architecture Behavioral of ROM_FC_84_81_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_81: ROM_ARRAY_PESOS_FC_84 := (
"10011110", 
"10010110", 
"10000110", 
"01111001", 
"01100111", 
"10011101", 
"10000111", 
"01111100", 
"01111110", 
"10100110", 
"01101011", 
"00101111", 
"10011011", 
"10001000", 
"10100111", 
"10000110", 
"10000010", 
"01111110", 
"01110101", 
"01110100", 
"01111010", 
"10001110", 
"10000010", 
"01010010", 
"10011000", 
"10010010", 
"10010011", 
"10011110", 
"01011100", 
"10110010", 
"10011010", 
"01110010", 
"01111001", 
"10010000", 
"10010010", 
"01111011", 
"01100110", 
"01011001", 
"10000010", 
"01111110", 
"10000100", 
"10101000", 
"10100110", 
"01010011", 
"10000111", 
"10100011", 
"01100001", 
"10010110", 
"01111010", 
"10001001", 
"01110010", 
"10001001", 
"10010111", 
"01100011", 
"01110100", 
"10000101", 
"01110101", 
"01101000", 
"10001001", 
"01110001", 
"01111110", 
"01110101", 
"10001110", 
"01011010", 
"10001101", 
"10000000", 
"10000000", 
"10011010", 
"10010101", 
"10000110", 
"01101101", 
"01101100", 
"01101110", 
"01100110", 
"10010111", 
"10011001", 
"01101100", 
"01110100", 
"10010001", 
"10000100", 
"01110000", 
"01001101", 
"01110000", 
"10100001", 
"00111011", 
"01011101", 
"10010100", 
"01101011", 
"10001000", 
"01000101", 
"01100110", 
"10000000", 
"01111110", 
"01100010", 
"01011101", 
"10001110", 
"01110100", 
"10001101", 
"10000000", 
"10011001", 
"01101000", 
"10100101", 
"01110010", 
"01101011", 
"01111101", 
"01110001", 
"01111011", 
"01110001", 
"01110011", 
"10010110", 
"01110100", 
"01101010", 
"01111101", 
"01110000", 
"01110010", 
"01110110", 
"01011001", 
"01010001", 
"01101111", 
"01011110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_81: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_81(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
