use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_31_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_31_LAYER;

architecture Behavioral of ROM_FC_120_31_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_31: ROM_ARRAY_PESOS_FC_120 := (
"01011000", 
"10001001", 
"10001001", 
"01111001", 
"01111011", 
"01011000", 
"01111011", 
"10000011", 
"01111110", 
"10001110", 
"10000000", 
"10001111", 
"10001000", 
"10000011", 
"01111011", 
"10000100", 
"01111000", 
"10010101", 
"01101011", 
"01001011", 
"10010001", 
"01100000", 
"10010000", 
"01011000", 
"01110111", 
"10001010", 
"10011001", 
"01110000", 
"10010001", 
"10011110", 
"01111101", 
"10000111", 
"01101000", 
"10011011", 
"10001011", 
"01101011", 
"10011010", 
"01100100", 
"10011111", 
"10001001", 
"01111111", 
"01101001", 
"01111001", 
"01100110", 
"01111011", 
"10011111", 
"10000011", 
"10010011", 
"01100001", 
"01101110", 
"10001111", 
"10000001", 
"01110011", 
"10001010", 
"01111100", 
"01110010", 
"01111110", 
"01000001", 
"10010001", 
"01001100", 
"01111001", 
"01111001", 
"10001001", 
"10011110", 
"01110001", 
"01101011", 
"01011110", 
"10100100", 
"10011000", 
"11000000", 
"10000100", 
"01100101", 
"01101100", 
"01110110", 
"10000111", 
"10000000", 
"01101111", 
"01101110", 
"10001011", 
"01101010", 
"10001110", 
"10100001", 
"01101111", 
"01101100", 
"10000001", 
"10000001", 
"01001001", 
"01111010", 
"10010011", 
"10100111", 
"01111000", 
"10010111", 
"01011000", 
"01111001", 
"10001100", 
"10000001", 
"01110100", 
"10111010", 
"10001110", 
"01010010", 
"01110000", 
"01010001", 
"10011001", 
"10000001", 
"10000100", 
"01010110", 
"01000001", 
"10011010", 
"01111001", 
"10001001", 
"10000101", 
"01110100", 
"01110010", 
"10010111", 
"00101101", 
"00111101", 
"10000010", 
"01111110", 
"10110111", 
"01010011", 
"01111001", 
"01111000", 
"01100100", 
"10101100", 
"00111000", 
"01011101", 
"10000011", 
"01101111", 
"10100010", 
"01001111", 
"01001000", 
"01110010", 
"01100000", 
"10010111", 
"10100110", 
"10001010", 
"10100110", 
"00101110", 
"10110010", 
"01001010", 
"10000011", 
"10000100", 
"01101111", 
"01101010", 
"10010010", 
"00111110", 
"10000101", 
"10000111", 
"10010011", 
"01110010", 
"10101010", 
"10001011", 
"10010110", 
"01010100", 
"01101000", 
"01101011", 
"01011101", 
"10011000", 
"01110111", 
"01101000", 
"10001110", 
"01100100", 
"01110101", 
"01010101", 
"01111110", 
"01111100", 
"10110101", 
"11101011", 
"01011010", 
"10001101", 
"00110110", 
"10011000", 
"01101010", 
"10011010", 
"01111101", 
"01101111", 
"10000110", 
"00011100", 
"01100010", 
"00110000", 
"01111111", 
"01111110", 
"10110000", 
"10110010", 
"01111100", 
"10001000", 
"01011001", 
"01011000", 
"01111011", 
"00111011", 
"10001100", 
"01110101", 
"01101010", 
"00010001", 
"11000000", 
"10010101", 
"10001000", 
"10100101", 
"01111010", 
"01011001", 
"10000011", 
"01011111", 
"10000010", 
"00011100", 
"10000010", 
"10001000", 
"10000101", 
"01011001", 
"01111101", 
"00110110", 
"10001110", 
"10011110", 
"01111111", 
"01110010", 
"01100111", 
"10010110", 
"10000101", 
"01110100", 
"01110111", 
"00111010", 
"10001110", 
"10111111", 
"01111110", 
"10010010", 
"01101010", 
"00001111", 
"10000110", 
"10011111", 
"01100110", 
"00101101", 
"10110011", 
"10101011", 
"01110000", 
"10001001", 
"00100100", 
"01001000", 
"10100011", 
"01011000", 
"01111110", 
"10001000", 
"10010001", 
"00101110", 
"11000111", 
"01100111", 
"01110011", 
"00011111", 
"00100101", 
"10011010", 
"01111011", 
"10010000", 
"01000011", 
"01111011", 
"01111111", 
"00111000", 
"01111011", 
"10001001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_31: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_31(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
