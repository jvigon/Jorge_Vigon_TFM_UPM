use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_28_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_28_LAYER;

architecture Behavioral of ROM_FC_84_28_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_28: ROM_ARRAY_PESOS_FC_84 := (
"01100101", 
"01111001", 
"01110100", 
"10000011", 
"01111000", 
"01110100", 
"10001001", 
"01110110", 
"10011111", 
"01110101", 
"01111010", 
"01111010", 
"01101011", 
"01101111", 
"01111001", 
"01111110", 
"01010000", 
"10010100", 
"01110001", 
"01011110", 
"01101001", 
"01011001", 
"01110011", 
"10001001", 
"01111001", 
"01110111", 
"01111110", 
"01101010", 
"01101000", 
"10001001", 
"10010011", 
"01101100", 
"01001111", 
"10001001", 
"01011001", 
"01001001", 
"10101000", 
"01101001", 
"10010010", 
"01101101", 
"01100001", 
"10110100", 
"01111001", 
"01110110", 
"10000111", 
"01001011", 
"10000100", 
"10000100", 
"01100011", 
"01100001", 
"10010111", 
"10000111", 
"01101100", 
"10010011", 
"01001011", 
"10100011", 
"01111000", 
"10001010", 
"01101101", 
"01110101", 
"01100001", 
"01100111", 
"01111010", 
"01001010", 
"01111010", 
"01011000", 
"10010001", 
"10011001", 
"10000010", 
"01111111", 
"01010100", 
"01100111", 
"01010101", 
"01100001", 
"10010010", 
"10010010", 
"01111110", 
"10001010", 
"01001101", 
"01111100", 
"01101000", 
"10000100", 
"01110000", 
"01100001", 
"01100100", 
"01111110", 
"10010110", 
"01010001", 
"10000111", 
"01001111", 
"01111000", 
"01110000", 
"01100111", 
"10011001", 
"01001111", 
"01101011", 
"01010111", 
"01110010", 
"01001100", 
"01100000", 
"10011000", 
"01101101", 
"01100100", 
"01110000", 
"01111111", 
"10010100", 
"01101111", 
"01101000", 
"01110101", 
"01101101", 
"01110010", 
"01100101", 
"01111000", 
"10001101", 
"10010011", 
"01101110", 
"01111100", 
"01111010", 
"10000111", 
"01011000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_28 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_28(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
