use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_96_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_96_LAYER;

architecture Behavioral of ROM_FC_120_96_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_96: ROM_ARRAY_PESOS_FC_120 := (
"10001111", 
"10001111", 
"01101101", 
"00110010", 
"10001111", 
"01110100", 
"01011110", 
"10000000", 
"10001100", 
"01101100", 
"10000011", 
"10100110", 
"10011110", 
"00111010", 
"01110110", 
"01101100", 
"10000011", 
"10000100", 
"10011101", 
"01111000", 
"10001111", 
"10000101", 
"01001010", 
"10001010", 
"01110011", 
"01101001", 
"01110000", 
"10101110", 
"01111111", 
"01011110", 
"10000011", 
"01110111", 
"01111010", 
"10111000", 
"10000001", 
"01101001", 
"01110101", 
"10010110", 
"01111001", 
"10000111", 
"10010000", 
"01001110", 
"10010011", 
"01010101", 
"10000100", 
"10101010", 
"10000100", 
"10001001", 
"10001110", 
"10010110", 
"01011010", 
"10100011", 
"10010010", 
"10000110", 
"01100110", 
"10001001", 
"10000100", 
"01001000", 
"10001110", 
"01110001", 
"01101000", 
"10101101", 
"10011010", 
"10110100", 
"01110111", 
"01111001", 
"01011010", 
"10111000", 
"10001111", 
"10000101", 
"01110000", 
"10000111", 
"10000010", 
"01010100", 
"01111010", 
"10001100", 
"10000110", 
"01110101", 
"10010100", 
"01101100", 
"01100100", 
"10011100", 
"01111110", 
"10001100", 
"10001001", 
"01110111", 
"01111000", 
"10000001", 
"10010001", 
"01110010", 
"01110110", 
"01110011", 
"10001000", 
"01010000", 
"01110010", 
"10001101", 
"10010010", 
"10011110", 
"01111000", 
"01111101", 
"10000001", 
"01110010", 
"01101100", 
"10000100", 
"10000011", 
"10001100", 
"10010111", 
"01011100", 
"10010010", 
"01010110", 
"10001011", 
"01111011", 
"01110111", 
"10001110", 
"01111101", 
"10001100", 
"01110111", 
"10010110", 
"10001101", 
"01111100", 
"10000101", 
"00110110", 
"01110100", 
"01000100", 
"01111110", 
"01101111", 
"10010010", 
"01111100", 
"01110011", 
"10001001", 
"01110000", 
"01111110", 
"10010010", 
"01111111", 
"10000001", 
"01011100", 
"10010010", 
"01101000", 
"01100000", 
"01111100", 
"01100111", 
"10000010", 
"01111011", 
"01110011", 
"01101100", 
"10000010", 
"01111110", 
"01110100", 
"10001111", 
"01011101", 
"01110110", 
"01101110", 
"10011000", 
"10000000", 
"01111100", 
"01101111", 
"10000010", 
"01100101", 
"10001101", 
"10001000", 
"01101111", 
"10010010", 
"10000011", 
"10100001", 
"01111100", 
"01100000", 
"10000011", 
"10001101", 
"01101111", 
"01011011", 
"01111010", 
"10001010", 
"10001010", 
"01100010", 
"10001001", 
"10000110", 
"01111110", 
"10000010", 
"01011001", 
"10011010", 
"10010101", 
"10100000", 
"01101100", 
"10011100", 
"10001010", 
"01010001", 
"01110111", 
"01100100", 
"01111110", 
"01111110", 
"10000010", 
"10000000", 
"01101110", 
"01111111", 
"10010100", 
"10000110", 
"01111100", 
"01100000", 
"00111000", 
"01101100", 
"01110001", 
"01010110", 
"10001001", 
"01010110", 
"01111010", 
"01111111", 
"01111010", 
"10010001", 
"10000010", 
"10011010", 
"10000100", 
"10010111", 
"10010011", 
"01010101", 
"10100001", 
"10010010", 
"01110100", 
"10000110", 
"01110011", 
"01110110", 
"01110101", 
"10000010", 
"01110010", 
"01110001", 
"10001001", 
"10010110", 
"10001100", 
"10000100", 
"01110111", 
"01010000", 
"10001010", 
"01100111", 
"01111101", 
"01110110", 
"01001010", 
"10111101", 
"10101010", 
"10100010", 
"01110110", 
"10001010", 
"10010001", 
"10101111", 
"01111011", 
"01001010", 
"10011000", 
"10001100", 
"01101011", 
"10010000", 
"01110110", 
"10011000", 
"01101100", 
"10100001", 
"10100110", 
"10010001", 
"01110100", 
"10000100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_96 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_96(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
