use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_29_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_29_LAYER;

architecture Behavioral of ROM_FC_84_29_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_29: ROM_ARRAY_PESOS_FC_84 := (
"10110110", 
"01110110", 
"01011110", 
"01110001", 
"10001011", 
"01111001", 
"01100111", 
"01100100", 
"01010000", 
"10101000", 
"10000001", 
"01111100", 
"01010100", 
"11000000", 
"01111011", 
"01100010", 
"10001101", 
"10000111", 
"10010010", 
"10000110", 
"01111111", 
"10000111", 
"01111000", 
"01010100", 
"10000111", 
"01110101", 
"01101011", 
"01101000", 
"10000011", 
"01100011", 
"10000110", 
"10000101", 
"01101101", 
"11010010", 
"01011111", 
"01010011", 
"01100010", 
"10010100", 
"01111001", 
"01110101", 
"01111100", 
"11000010", 
"01111101", 
"01001110", 
"01001010", 
"01010001", 
"10010100", 
"01101010", 
"01100110", 
"10001101", 
"01101001", 
"01111101", 
"01101011", 
"01010100", 
"10000110", 
"10011011", 
"01101110", 
"01111110", 
"01010000", 
"11001100", 
"10001000", 
"01100100", 
"10000110", 
"01011000", 
"10010011", 
"00101010", 
"10110001", 
"10010000", 
"10001000", 
"10000010", 
"10000111", 
"10011010", 
"01011000", 
"10000000", 
"10011101", 
"01111001", 
"01111100", 
"10110011", 
"01011110", 
"10000111", 
"01101000", 
"10001011", 
"01111010", 
"01110101", 
"10010011", 
"10001001", 
"01110110", 
"10010101", 
"01111101", 
"10001101", 
"01111010", 
"11011110", 
"10010101", 
"01110100", 
"01000110", 
"10000011", 
"10000100", 
"01101001", 
"01000101", 
"01100011", 
"10011011", 
"01111101", 
"01100011", 
"01011110", 
"01100001", 
"01101110", 
"01101100", 
"10010001", 
"10011000", 
"10011001", 
"10000011", 
"01100010", 
"01101100", 
"00010110", 
"10010110", 
"10000110", 
"01001001", 
"01100011", 
"10011010", 
"10001011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_29 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_29(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
