use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_18_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_18_LAYER;

architecture Behavioral of ROM_FC_120_18_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_18: ROM_ARRAY_PESOS_FC_120 := (
"01111110", 
"10011010", 
"01100001", 
"01100011", 
"01100011", 
"10011001", 
"01101001", 
"11001000", 
"01111110", 
"01110101", 
"01101001", 
"01000111", 
"01110100", 
"01001110", 
"01101110", 
"01111101", 
"01100111", 
"01011100", 
"01011110", 
"00111101", 
"01101000", 
"01011111", 
"10011000", 
"10011100", 
"10001001", 
"01101110", 
"00111011", 
"00111010", 
"01010001", 
"01101011", 
"01101110", 
"10001011", 
"10100101", 
"01111001", 
"01000011", 
"01100000", 
"10100101", 
"01111100", 
"10001010", 
"01010011", 
"01101100", 
"01100000", 
"10000001", 
"01101111", 
"01110110", 
"01100000", 
"01101011", 
"10010001", 
"10000011", 
"00111110", 
"01111001", 
"01101100", 
"10001000", 
"10000000", 
"01110101", 
"10100100", 
"10001111", 
"10001111", 
"10001001", 
"01110011", 
"10001000", 
"10010001", 
"10000001", 
"10011011", 
"01010001", 
"01110001", 
"10001010", 
"01100101", 
"10101000", 
"01011011", 
"10100111", 
"10110001", 
"01101110", 
"01111011", 
"01011110", 
"01000000", 
"10010100", 
"01010010", 
"10010111", 
"01110111", 
"10110100", 
"10011100", 
"01100010", 
"01010011", 
"11000001", 
"10010110", 
"10001010", 
"10010111", 
"01011111", 
"10001111", 
"01100011", 
"01111010", 
"01100001", 
"00110001", 
"01111010", 
"10001111", 
"10100101", 
"10010000", 
"01101010", 
"10100110", 
"01111110", 
"10000011", 
"10101011", 
"10010101", 
"10010101", 
"01111111", 
"10000101", 
"10000010", 
"01010100", 
"01101101", 
"01110100", 
"01101010", 
"10001011", 
"01110101", 
"10001110", 
"10101000", 
"10000000", 
"01110111", 
"10010110", 
"01010000", 
"10001110", 
"01011101", 
"01010011", 
"10100011", 
"10000110", 
"10110010", 
"10001011", 
"01110111", 
"10010100", 
"01110111", 
"01001111", 
"10011001", 
"10100101", 
"01110000", 
"01110100", 
"01110010", 
"01111101", 
"10011001", 
"01110000", 
"01011100", 
"01011110", 
"10011100", 
"01011011", 
"01110011", 
"01100010", 
"01100110", 
"01111101", 
"10010100", 
"10000100", 
"01011010", 
"01011111", 
"10100110", 
"10010001", 
"01110111", 
"01110110", 
"01101100", 
"01101101", 
"01010011", 
"10001110", 
"10010011", 
"01100010", 
"10000010", 
"10010001", 
"01110011", 
"10001110", 
"10000001", 
"01100100", 
"01010001", 
"10000010", 
"10000110", 
"01101011", 
"01101101", 
"10110111", 
"10001001", 
"10100011", 
"10010100", 
"10011110", 
"10001110", 
"10001011", 
"01100111", 
"01110000", 
"01100001", 
"10001000", 
"01111111", 
"10000011", 
"10100010", 
"10001110", 
"10100011", 
"11000110", 
"10001001", 
"10000010", 
"10001000", 
"10001111", 
"10000100", 
"01111011", 
"11000111", 
"01110011", 
"01010101", 
"01101010", 
"01010110", 
"10001010", 
"10000000", 
"10000101", 
"01111110", 
"10000011", 
"10010011", 
"01111001", 
"10000100", 
"01100101", 
"01011010", 
"10011011", 
"10011001", 
"10001100", 
"01100000", 
"01011001", 
"00111000", 
"10000010", 
"10011101", 
"10010111", 
"10011000", 
"10101011", 
"10000101", 
"01110110", 
"01111000", 
"10011000", 
"10010101", 
"10011100", 
"01001011", 
"01100100", 
"10100001", 
"01010010", 
"10110000", 
"10110111", 
"10011011", 
"10010111", 
"10000111", 
"10000001", 
"01001111", 
"01110010", 
"10000010", 
"01011111", 
"10010100", 
"01100100", 
"10000011", 
"01111001", 
"01100011", 
"01000010", 
"11001101", 
"01111010", 
"01011010", 
"10010001", 
"10011101", 
"01010111", 
"01000010", 
"10001011", 
"01110001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_18: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_18(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
