use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_34_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_34_LAYER;

architecture Behavioral of ROM_FC_84_34_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_34: ROM_ARRAY_PESOS_FC_84 := (
"10101010", 
"01110010", 
"01111011", 
"01110101", 
"01110111", 
"01110111", 
"10001000", 
"01100101", 
"01111011", 
"11101100", 
"01110011", 
"01111001", 
"10011011", 
"01100111", 
"01011010", 
"10101111", 
"01111110", 
"01101110", 
"01101010", 
"10000001", 
"10110010", 
"01011000", 
"10111110", 
"01011001", 
"10010010", 
"10010110", 
"10000111", 
"10000010", 
"01010101", 
"10100001", 
"10011000", 
"00111011", 
"01100110", 
"10000110", 
"10000101", 
"10000011", 
"10111000", 
"10000010", 
"10000000", 
"10001100", 
"10010101", 
"10010101", 
"01010100", 
"01101101", 
"10100101", 
"10000101", 
"01110001", 
"10001011", 
"01010000", 
"01111110", 
"01001001", 
"01100110", 
"01111001", 
"10001000", 
"01101100", 
"01110100", 
"10000110", 
"01101110", 
"01101100", 
"10010001", 
"01011010", 
"01101011", 
"01111111", 
"01001011", 
"01001111", 
"10001010", 
"01111111", 
"10001111", 
"10011110", 
"10111001", 
"01111010", 
"00111101", 
"10000110", 
"01110101", 
"01110010", 
"10011000", 
"10101111", 
"10000110", 
"10010000", 
"01110001", 
"10010100", 
"10001111", 
"10101011", 
"10010011", 
"01101101", 
"10000010", 
"10010010", 
"01101111", 
"10000110", 
"01101001", 
"01111101", 
"01000111", 
"10111010", 
"01000101", 
"01011001", 
"01110100", 
"01111101", 
"10001001", 
"10010000", 
"10110110", 
"01101011", 
"01111101", 
"10011111", 
"10001011", 
"01001001", 
"10000111", 
"01110101", 
"10000011", 
"10001000", 
"01100000", 
"10001000", 
"10000011", 
"01111100", 
"01111111", 
"10011111", 
"01100001", 
"10100110", 
"01101100", 
"01101010", 
"01110111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_34 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_34(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
