use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_82_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_82_LAYER;

architecture Behavioral of ROM_FC_120_82_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_82: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"01111001", 
"01100011", 
"01101011", 
"10001110", 
"01000011", 
"01110000", 
"01101111", 
"01101100", 
"10001001", 
"10011100", 
"11001110", 
"01111111", 
"01100101", 
"10000010", 
"10010010", 
"01111100", 
"10001100", 
"01011110", 
"01111101", 
"10100010", 
"10001000", 
"01110001", 
"01100010", 
"10010001", 
"10000011", 
"10001010", 
"10100001", 
"10010011", 
"01011001", 
"01101010", 
"01111011", 
"01111000", 
"10010011", 
"10000111", 
"10100010", 
"10010001", 
"10001111", 
"01011000", 
"01111110", 
"10000101", 
"10011010", 
"01110001", 
"10110000", 
"01101111", 
"11001101", 
"10011010", 
"01110111", 
"10000111", 
"10011000", 
"01110111", 
"01010101", 
"01111111", 
"10011011", 
"01011011", 
"01110101", 
"01110000", 
"01100101", 
"01100111", 
"01101101", 
"01101011", 
"10101110", 
"10010011", 
"10011000", 
"10001110", 
"10000010", 
"01111101", 
"01111010", 
"01100011", 
"01100111", 
"10010011", 
"10110001", 
"10000110", 
"01100100", 
"01110100", 
"01110001", 
"10000100", 
"10000101", 
"01110110", 
"10000000", 
"01100101", 
"10000001", 
"01101111", 
"01111101", 
"01100101", 
"10000010", 
"01111001", 
"10000011", 
"10001000", 
"01101111", 
"01110111", 
"01010101", 
"01101100", 
"10011101", 
"01111111", 
"10000001", 
"10011000", 
"01111010", 
"01100000", 
"01101011", 
"01110011", 
"01110110", 
"10001011", 
"10010000", 
"01111000", 
"01111011", 
"01110110", 
"01110000", 
"10001010", 
"11000001", 
"01110000", 
"01100101", 
"10100001", 
"10000001", 
"01101010", 
"01011100", 
"01101110", 
"10000010", 
"10100010", 
"10001011", 
"10000000", 
"01111010", 
"01110000", 
"01101111", 
"01101001", 
"01101111", 
"01101100", 
"01101110", 
"01101000", 
"10000111", 
"01110101", 
"01110011", 
"10110100", 
"01010101", 
"11000111", 
"10110011", 
"01101110", 
"10000100", 
"10000101", 
"10010110", 
"10110010", 
"01011000", 
"10000101", 
"01111001", 
"10011110", 
"10110101", 
"10010110", 
"10000001", 
"01110001", 
"01101101", 
"01110111", 
"10001011", 
"01101000", 
"10011100", 
"01110011", 
"01110011", 
"10001101", 
"00111100", 
"10000011", 
"10000010", 
"10010100", 
"10000100", 
"01111110", 
"01111111", 
"10010000", 
"10000100", 
"01100010", 
"10010101", 
"10010001", 
"01110000", 
"10000011", 
"01100011", 
"01111110", 
"01100001", 
"01110101", 
"01111100", 
"10000110", 
"01001101", 
"01110010", 
"11000100", 
"10001110", 
"01110011", 
"01110111", 
"10011000", 
"10000111", 
"10000000", 
"01111101", 
"01101101", 
"01101111", 
"01011101", 
"01110111", 
"10001100", 
"01100011", 
"10001000", 
"01101011", 
"10011001", 
"01101100", 
"10001000", 
"01111011", 
"10010110", 
"10010000", 
"10000000", 
"10010010", 
"01111101", 
"01011101", 
"01110011", 
"01110010", 
"01101101", 
"10011101", 
"10011110", 
"01110101", 
"10000100", 
"01111001", 
"10010100", 
"01111101", 
"10011001", 
"01100000", 
"10000000", 
"01111110", 
"01110010", 
"01101011", 
"10000001", 
"01111111", 
"01111010", 
"01100011", 
"10000101", 
"01101110", 
"01111101", 
"10000110", 
"10000000", 
"01110100", 
"01110111", 
"10010111", 
"01111100", 
"10001000", 
"01100000", 
"01110010", 
"01101101", 
"10001000", 
"10000000", 
"00110001", 
"00101111", 
"10100011", 
"11010111", 
"01101100", 
"01110011", 
"01011100", 
"01011001", 
"10000110", 
"11000001", 
"10001110", 
"10000111", 
"01111100", 
"10001101", 
"01111001", 
"01111000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_82: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_82(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
