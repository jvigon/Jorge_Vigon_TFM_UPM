use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_1_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_1_LAYER;

architecture Behavioral of ROM_FC_120_1_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_1: ROM_ARRAY_PESOS_FC_120 := (
"10010111", 
"10011010", 
"01011011", 
"01100100", 
"10100010", 
"11010001", 
"01110100", 
"01110111", 
"10001000", 
"10000011", 
"10101001", 
"10011001", 
"01101000", 
"01100000", 
"10000110", 
"10011010", 
"01111111", 
"10001011", 
"01100010", 
"01110111", 
"01001101", 
"10110111", 
"01110111", 
"01100001", 
"10000101", 
"01011100", 
"01010001", 
"10111000", 
"01011100", 
"10111010", 
"10100101", 
"10001000", 
"10111011", 
"10001010", 
"01110010", 
"10110101", 
"01101100", 
"10000110", 
"10111001", 
"10001100", 
"10001000", 
"01100001", 
"01101101", 
"01110100", 
"01011100", 
"01011111", 
"01110000", 
"01110100", 
"10011111", 
"10010101", 
"01101010", 
"10100000", 
"10101101", 
"01100000", 
"11000011", 
"10100111", 
"01101000", 
"10010111", 
"01110001", 
"01110100", 
"10001000", 
"01101111", 
"01111000", 
"10000010", 
"01110010", 
"10111000", 
"01110101", 
"10011000", 
"10000101", 
"01111011", 
"10011110", 
"01100100", 
"01100101", 
"01100000", 
"10101001", 
"11000011", 
"10001101", 
"01010001", 
"01111111", 
"10001011", 
"01100000", 
"10010101", 
"10001011", 
"10001111", 
"10001110", 
"01101100", 
"10001111", 
"01111100", 
"01101110", 
"01100001", 
"01110101", 
"10100010", 
"10100001", 
"01110000", 
"01110000", 
"01101101", 
"01100101", 
"01011111", 
"01111100", 
"10000011", 
"10010101", 
"01011110", 
"01100011", 
"01111010", 
"10010101", 
"10011000", 
"10001011", 
"01110011", 
"01110101", 
"01001011", 
"01110111", 
"10001010", 
"01110000", 
"00111010", 
"10100110", 
"10011010", 
"10011111", 
"01001101", 
"01100100", 
"10000111", 
"01111011", 
"10011100", 
"01110011", 
"01101110", 
"00111001", 
"01011110", 
"01101101", 
"10001100", 
"01011101", 
"10001001", 
"01011100", 
"01101011", 
"10111010", 
"10000001", 
"10101001", 
"01001010", 
"01100001", 
"10100010", 
"10000111", 
"10110000", 
"01101011", 
"01011000", 
"10010010", 
"01110111", 
"01010001", 
"10001101", 
"10011111", 
"10011111", 
"10001000", 
"01100110", 
"01101100", 
"01100110", 
"01110110", 
"01101110", 
"10001010", 
"01111101", 
"01100110", 
"00011101", 
"10001101", 
"10000110", 
"01100100", 
"10011101", 
"10000100", 
"01110011", 
"01110100", 
"01100111", 
"10000011", 
"10010001", 
"10001100", 
"10010100", 
"10101100", 
"10000001", 
"01111111", 
"01111000", 
"01101000", 
"10000011", 
"01101010", 
"01111000", 
"01111000", 
"01111010", 
"01111110", 
"01010101", 
"01110101", 
"10001111", 
"01110001", 
"10100110", 
"10000000", 
"01101010", 
"10000101", 
"10010000", 
"10011101", 
"10000001", 
"01011101", 
"01110101", 
"01011110", 
"01011010", 
"10000001", 
"00100110", 
"10100000", 
"10000011", 
"01110111", 
"10001011", 
"01110000", 
"10000101", 
"01000010", 
"10000010", 
"10011010", 
"01111011", 
"01110101", 
"01110111", 
"01101001", 
"10100000", 
"01111101", 
"01111101", 
"10011001", 
"01001100", 
"10000100", 
"01110001", 
"10001011", 
"01111001", 
"01011001", 
"10011000", 
"10000101", 
"01111100", 
"10110001", 
"01111101", 
"10101000", 
"10000110", 
"01111100", 
"10010010", 
"01111100", 
"10001100", 
"10000001", 
"01101011", 
"10001111", 
"01110010", 
"01101000", 
"01101001", 
"10000011", 
"10010100", 
"10000110", 
"10011011", 
"10000010", 
"01001000", 
"01110111", 
"01111011", 
"10000011", 
"10000010", 
"01101110", 
"10011001", 
"01100100", 
"10010011", 
"10101110", 
"10011101", 
"01101111", 
"01111111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_1 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_1(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
