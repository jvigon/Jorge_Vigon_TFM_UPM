use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_38_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_38_LAYER;

architecture Behavioral of ROM_FC_84_38_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_38: ROM_ARRAY_PESOS_FC_84 := (
"01101101", 
"01100110", 
"10000111", 
"10000010", 
"10001001", 
"10001011", 
"01101000", 
"01001111", 
"01011111", 
"01110010", 
"10010000", 
"10110101", 
"01011011", 
"01011011", 
"01110001", 
"01111010", 
"01111011", 
"10011011", 
"00111010", 
"10001111", 
"01101011", 
"01100000", 
"10001100", 
"01101010", 
"01101110", 
"01100111", 
"01011000", 
"01101110", 
"01100110", 
"01100111", 
"01100011", 
"10011110", 
"10000111", 
"01110000", 
"01110011", 
"01001100", 
"01100010", 
"01101001", 
"10110011", 
"10010000", 
"01001000", 
"01110111", 
"10010110", 
"01001111", 
"01011100", 
"10000000", 
"01011010", 
"10001011", 
"01000000", 
"01111011", 
"01110111", 
"10000011", 
"10000101", 
"01111110", 
"01101111", 
"01100110", 
"01100100", 
"10010111", 
"10000110", 
"10000000", 
"01101111", 
"01110000", 
"10010010", 
"01111000", 
"01010110", 
"01001110", 
"10000011", 
"10010110", 
"01111000", 
"01110000", 
"01101010", 
"01101010", 
"01101000", 
"10010011", 
"10001100", 
"01110111", 
"01100010", 
"10010010", 
"10001100", 
"01011100", 
"10000011", 
"10001101", 
"01010010", 
"01110000", 
"01001111", 
"01011111", 
"10000110", 
"10011011", 
"10001111", 
"01100011", 
"10001001", 
"10000111", 
"10010011", 
"01010110", 
"01011110", 
"01110101", 
"01011000", 
"01110011", 
"10011001", 
"01110010", 
"01101100", 
"01101110", 
"10101011", 
"01110111", 
"10000000", 
"10010011", 
"01101101", 
"01111101", 
"10010110", 
"10000011", 
"01110001", 
"01111011", 
"10001111", 
"10010001", 
"10001100", 
"01011111", 
"01010111", 
"10001000", 
"10001101", 
"01100111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_38: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_38(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
