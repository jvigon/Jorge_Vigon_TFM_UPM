use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_48_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_48_LAYER;

architecture Behavioral of ROM_FC_84_48_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_48: ROM_ARRAY_PESOS_FC_84 := (
"01011000", 
"10010100", 
"01110001", 
"10000010", 
"01100110", 
"01110110", 
"10001010", 
"01010001", 
"01100110", 
"01101000", 
"01110110", 
"01101000", 
"01110111", 
"10001010", 
"01110100", 
"01100110", 
"10000111", 
"10000011", 
"01101110", 
"10010010", 
"01101010", 
"10101101", 
"10000110", 
"01001101", 
"10001101", 
"01101100", 
"10000001", 
"01101010", 
"01111001", 
"10000101", 
"01101110", 
"01110111", 
"10001001", 
"10010011", 
"10011101", 
"01100011", 
"10001000", 
"10000111", 
"01100100", 
"01101101", 
"01011110", 
"10000111", 
"10010010", 
"10000010", 
"01011110", 
"01001111", 
"10001000", 
"10000100", 
"10000101", 
"10000011", 
"01111000", 
"01101010", 
"10000011", 
"01011111", 
"01001001", 
"01010100", 
"01110001", 
"10010011", 
"01110110", 
"10011000", 
"10001001", 
"01101100", 
"01110010", 
"01011001", 
"01101000", 
"01000111", 
"01100110", 
"10000001", 
"01110000", 
"01111011", 
"01111100", 
"01010100", 
"10000100", 
"01101110", 
"01110001", 
"01110001", 
"01110000", 
"01110110", 
"01110001", 
"01101110", 
"10010000", 
"01001010", 
"01010111", 
"01011111", 
"01010101", 
"01011101", 
"01111000", 
"01100010", 
"01101111", 
"01110111", 
"01010110", 
"01101010", 
"01101010", 
"01110010", 
"10001010", 
"10010101", 
"01110010", 
"01101110", 
"01100111", 
"01101110", 
"01101101", 
"01110000", 
"01010001", 
"01100100", 
"01111010", 
"01100001", 
"10000010", 
"01111001", 
"01100111", 
"10001000", 
"01100010", 
"10000010", 
"01110101", 
"01110000", 
"10011101", 
"10000011", 
"01001100", 
"10011010", 
"10001110", 
"01011101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_48: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_48(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
