use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_80_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_80_LAYER;

architecture Behavioral of ROM_FC_120_80_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_80: ROM_ARRAY_PESOS_FC_120 := (
"01111001", 
"01110011", 
"10011111", 
"10101010", 
"01111111", 
"01100110", 
"01100000", 
"01110010", 
"01110001", 
"01010011", 
"01101110", 
"10111110", 
"10011011", 
"01111111", 
"01101011", 
"01101001", 
"01110101", 
"01110011", 
"01110100", 
"01111000", 
"01111000", 
"10001000", 
"01110001", 
"01110110", 
"10000100", 
"01101101", 
"01100011", 
"10001100", 
"01110010", 
"01111001", 
"01110101", 
"01110000", 
"10001111", 
"01101010", 
"00110111", 
"01101110", 
"01101111", 
"10000100", 
"01100100", 
"01111001", 
"01111011", 
"01011010", 
"01001110", 
"01011000", 
"01110110", 
"10001100", 
"01111000", 
"10001010", 
"01100111", 
"01101001", 
"01101011", 
"01111111", 
"01101001", 
"01111011", 
"01110110", 
"10001010", 
"01110010", 
"01001000", 
"01110000", 
"01110010", 
"00111000", 
"10000100", 
"01110011", 
"10001001", 
"01111111", 
"01111011", 
"10011110", 
"10001101", 
"01110010", 
"01100111", 
"01100000", 
"10001101", 
"01110010", 
"01111101", 
"10001001", 
"01110010", 
"10000111", 
"10000110", 
"01110001", 
"01110000", 
"01111101", 
"01100111", 
"01111000", 
"10000000", 
"10001001", 
"01101001", 
"01010100", 
"10000100", 
"10001111", 
"01100111", 
"01011111", 
"01101101", 
"01101010", 
"01010111", 
"10000000", 
"01111001", 
"10000011", 
"01011011", 
"01100111", 
"01100010", 
"10001101", 
"01010111", 
"01011111", 
"10000100", 
"10010000", 
"10001011", 
"01101011", 
"01110011", 
"01110100", 
"01100101", 
"10000010", 
"10001111", 
"01100110", 
"01001100", 
"01101101", 
"10011000", 
"01110101", 
"01010010", 
"10000010", 
"01110100", 
"01101001", 
"00110101", 
"01011001", 
"01110100", 
"10001001", 
"01110111", 
"01101000", 
"10000000", 
"01110001", 
"01100110", 
"01010110", 
"01100100", 
"10000000", 
"01110011", 
"10010000", 
"10001101", 
"01110010", 
"10000100", 
"01100111", 
"10110101", 
"10010100", 
"01101001", 
"10001011", 
"01111001", 
"01111010", 
"01100111", 
"01010100", 
"01010010", 
"01110010", 
"10000011", 
"01101011", 
"01111010", 
"10001011", 
"01010011", 
"01001011", 
"10000001", 
"10010011", 
"01111101", 
"01100011", 
"01111111", 
"10000001", 
"10001110", 
"01011001", 
"01011001", 
"01111001", 
"01111100", 
"01100010", 
"01011011", 
"01111100", 
"01010110", 
"01110100", 
"01101101", 
"10000100", 
"01101110", 
"01111010", 
"01101100", 
"10000001", 
"10001111", 
"10000010", 
"00100100", 
"01111101", 
"01101100", 
"01100011", 
"01110101", 
"10001110", 
"01110000", 
"01100000", 
"01100110", 
"10100111", 
"00111110", 
"01101011", 
"10001100", 
"10001010", 
"01110011", 
"01111111", 
"01001100", 
"10010010", 
"10000100", 
"10000110", 
"01101010", 
"01101001", 
"01110100", 
"01011101", 
"01110100", 
"10011111", 
"10101110", 
"10000010", 
"01111011", 
"10000011", 
"10001000", 
"10110000", 
"01111100", 
"01110110", 
"01101100", 
"01011100", 
"01100001", 
"10000101", 
"10010001", 
"01111000", 
"01011111", 
"10011000", 
"01100011", 
"01111100", 
"10000110", 
"10000101", 
"10001001", 
"01111001", 
"01111101", 
"10001010", 
"01100001", 
"01101010", 
"01100011", 
"01111001", 
"10000000", 
"01110010", 
"01000110", 
"10110010", 
"10001100", 
"01111110", 
"01110010", 
"01110100", 
"01100001", 
"10100110", 
"10001000", 
"10000100", 
"01110011", 
"01100010", 
"01110101", 
"01110000", 
"10010010", 
"01111100", 
"00111011", 
"11000011", 
"10001010", 
"01101110", 
"01110111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_80: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_80(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
