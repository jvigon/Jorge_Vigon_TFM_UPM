use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_38_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_38_LAYER;

architecture Behavioral of ROM_FC_120_38_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_38: ROM_ARRAY_PESOS_FC_120 := (
"10010100", 
"10001011", 
"01101100", 
"10010100", 
"01010001", 
"01111101", 
"01110011", 
"01101010", 
"10001010", 
"10010100", 
"01101011", 
"10101010", 
"01011101", 
"11011100", 
"01110010", 
"10010011", 
"10000100", 
"10101100", 
"01011101", 
"01010110", 
"01101001", 
"01110010", 
"10010101", 
"10000001", 
"01100111", 
"10001100", 
"01101110", 
"10100000", 
"10000111", 
"01110001", 
"10001101", 
"10000000", 
"10000100", 
"10000110", 
"01000011", 
"00111010", 
"01100010", 
"01111100", 
"10011101", 
"01011101", 
"01110111", 
"01110000", 
"01010001", 
"10011011", 
"10100101", 
"01011001", 
"10011001", 
"01100101", 
"10001100", 
"10001011", 
"01101110", 
"01010000", 
"01110011", 
"10111001", 
"01111100", 
"01101100", 
"01111010", 
"10000011", 
"01110010", 
"01011101", 
"10001100", 
"01010111", 
"01010111", 
"10010000", 
"01101110", 
"10011110", 
"01101100", 
"01100011", 
"01001101", 
"01011110", 
"10010100", 
"10001101", 
"01111111", 
"01111110", 
"10000101", 
"10000110", 
"10000010", 
"01111011", 
"10001100", 
"01101101", 
"01100100", 
"01110100", 
"01010011", 
"00110101", 
"01110011", 
"10011000", 
"10001110", 
"01110100", 
"01100101", 
"01101110", 
"10010100", 
"10011100", 
"10000001", 
"01110101", 
"01111110", 
"01110011", 
"10100100", 
"10000111", 
"01110010", 
"00011011", 
"01110110", 
"10000010", 
"10000001", 
"01101010", 
"01101110", 
"10010001", 
"10011010", 
"10010010", 
"01111101", 
"01011110", 
"01111011", 
"01111111", 
"10001110", 
"10100101", 
"01110000", 
"01011111", 
"01011111", 
"01110000", 
"01111100", 
"10001010", 
"01111110", 
"01111011", 
"10100111", 
"10001101", 
"10001010", 
"00110010", 
"10001000", 
"01101100", 
"01101111", 
"01110101", 
"01000011", 
"01010011", 
"10011011", 
"10001110", 
"10010100", 
"10100001", 
"10111011", 
"10001110", 
"01001101", 
"01101111", 
"01111100", 
"10001110", 
"10001100", 
"01101010", 
"11010101", 
"10001100", 
"01111111", 
"01011100", 
"01101111", 
"10000101", 
"01111100", 
"10011010", 
"01010110", 
"10000100", 
"10001001", 
"01101110", 
"01101101", 
"10011001", 
"10000101", 
"01111001", 
"10110001", 
"01101001", 
"01101111", 
"01011010", 
"10001001", 
"10000110", 
"01010111", 
"10001000", 
"10000110", 
"10000010", 
"01111010", 
"01100100", 
"10000000", 
"00100111", 
"01111001", 
"01101100", 
"10010000", 
"01000100", 
"01111011", 
"01110010", 
"01110011", 
"01101110", 
"10011110", 
"10000101", 
"01101101", 
"01101000", 
"10000010", 
"01111111", 
"10010110", 
"01011110", 
"01110100", 
"01101111", 
"01111110", 
"01110101", 
"01100001", 
"01111011", 
"01101110", 
"10110001", 
"10011100", 
"10111010", 
"10100101", 
"01100101", 
"01110011", 
"01111101", 
"01011100", 
"01100101", 
"01110010", 
"10001110", 
"11000010", 
"01100101", 
"00011110", 
"01110100", 
"01010111", 
"10011111", 
"01111111", 
"10111100", 
"01101001", 
"01101100", 
"10011101", 
"01100001", 
"00111011", 
"01010111", 
"10000000", 
"10000110", 
"01101100", 
"00010111", 
"01010101", 
"01010001", 
"01100110", 
"10000001", 
"01101110", 
"01111111", 
"10011101", 
"01101111", 
"10000011", 
"01010001", 
"01110100", 
"10011001", 
"01111001", 
"10000111", 
"00111011", 
"00101010", 
"10001011", 
"01111010", 
"01111001", 
"00110000", 
"10100100", 
"01011000", 
"01110001", 
"01111111", 
"01011000", 
"10101000", 
"01110111", 
"01100000", 
"10001110", 
"01101010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_38: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_38(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
