use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_66_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_66_LAYER;

architecture Behavioral of ROM_FC_84_66_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_66: ROM_ARRAY_PESOS_FC_84 := (
"01000110", 
"01111000", 
"10100000", 
"01111100", 
"01100010", 
"01111001", 
"01110010", 
"01110111", 
"10011010", 
"01110100", 
"10100111", 
"01010001", 
"01001101", 
"10001011", 
"01101001", 
"10000000", 
"01010101", 
"10011100", 
"10000110", 
"01010011", 
"01111110", 
"10001001", 
"01101100", 
"01101001", 
"01111110", 
"10100101", 
"01011001", 
"01111000", 
"01010000", 
"10011011", 
"10111011", 
"01011100", 
"01000010", 
"10001101", 
"01100110", 
"01011010", 
"01100110", 
"01110001", 
"01111001", 
"01001101", 
"01001110", 
"10010111", 
"01010001", 
"10001110", 
"01001100", 
"01101010", 
"01101011", 
"10010110", 
"10000111", 
"01110111", 
"01100010", 
"10000100", 
"01111111", 
"01111111", 
"10001001", 
"10001100", 
"01110110", 
"10000000", 
"01001011", 
"10011111", 
"10000000", 
"10001000", 
"01100011", 
"01000011", 
"10011000", 
"01011001", 
"10011101", 
"01100010", 
"10011001", 
"01110100", 
"01100101", 
"01110000", 
"10011111", 
"01000011", 
"01010000", 
"01101110", 
"01011111", 
"10000110", 
"10011001", 
"01011111", 
"01010101", 
"01101110", 
"01110110", 
"01101111", 
"01110011", 
"01101110", 
"01111111", 
"10000101", 
"10010000", 
"10000100", 
"01100110", 
"11001000", 
"10001010", 
"10010010", 
"01111000", 
"01110100", 
"10000111", 
"10001011", 
"01100100", 
"01111100", 
"10010011", 
"10001100", 
"01010101", 
"01000111", 
"10001000", 
"01011010", 
"01111010", 
"01010001", 
"01011110", 
"01101111", 
"01011010", 
"01011010", 
"01101111", 
"10010100", 
"10000110", 
"01111010", 
"10001101", 
"10011100", 
"10010110", 
"10000010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_66: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_66(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
