use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_84_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_84_LAYER;

architecture Behavioral of ROM_FC_120_84_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_84: ROM_ARRAY_PESOS_FC_120 := (
"01111100", 
"01100001", 
"01100111", 
"01100101", 
"01111010", 
"01010111", 
"10011000", 
"10000001", 
"01111011", 
"01111000", 
"01101110", 
"01101111", 
"10001011", 
"00101111", 
"10000100", 
"01111001", 
"01111111", 
"01110100", 
"10010000", 
"01110100", 
"10000001", 
"01010110", 
"10000100", 
"10100111", 
"10001101", 
"10010001", 
"10111001", 
"01010101", 
"10100010", 
"00011000", 
"01110010", 
"01100100", 
"01011000", 
"01011010", 
"10011000", 
"01111111", 
"01110000", 
"01001010", 
"00110100", 
"01111000", 
"10010110", 
"10101101", 
"10001111", 
"01100101", 
"10001001", 
"10000001", 
"10000010", 
"10001110", 
"01001011", 
"01010110", 
"10000010", 
"10000100", 
"10001010", 
"00110110", 
"00001011", 
"10011000", 
"10010101", 
"10011101", 
"01110000", 
"10000001", 
"01000111", 
"10001001", 
"10001101", 
"01111001", 
"10000101", 
"01000001", 
"01111010", 
"01111010", 
"01110111", 
"10100010", 
"01110000", 
"01011011", 
"10010111", 
"10000100", 
"10000100", 
"01011110", 
"00011101", 
"10010011", 
"10000110", 
"01110000", 
"10000110", 
"01101110", 
"10000011", 
"10101110", 
"10000110", 
"01111111", 
"01111100", 
"01101001", 
"10010001", 
"10100011", 
"10001100", 
"01101111", 
"01010111", 
"01100010", 
"01110010", 
"01101010", 
"10010010", 
"10000001", 
"01111010", 
"10000111", 
"01100111", 
"01110001", 
"01001001", 
"10001110", 
"01110110", 
"01111001", 
"10001011", 
"10001000", 
"01110010", 
"10000010", 
"01111101", 
"01110010", 
"01110001", 
"10010010", 
"01011100", 
"01010110", 
"01101100", 
"10000111", 
"10010111", 
"01101010", 
"10010010", 
"10010101", 
"01010010", 
"10100011", 
"10010011", 
"10010010", 
"10000010", 
"01111000", 
"01100000", 
"01101001", 
"10101011", 
"01111011", 
"01111001", 
"01110110", 
"01000010", 
"01011101", 
"10001111", 
"10000100", 
"10000011", 
"01111110", 
"01010110", 
"01110000", 
"01110001", 
"10010000", 
"01111001", 
"01010011", 
"01111010", 
"10011011", 
"01110011", 
"10011101", 
"01110001", 
"01111001", 
"10001100", 
"10100010", 
"01010110", 
"10000001", 
"01101100", 
"10000111", 
"01110101", 
"10000101", 
"01110100", 
"10010101", 
"10000010", 
"10001001", 
"01100111", 
"10001000", 
"01110101", 
"01111010", 
"10001101", 
"01100100", 
"01110111", 
"10000010", 
"10000101", 
"10100001", 
"10000100", 
"01101101", 
"01111100", 
"10011100", 
"01110011", 
"01000111", 
"10001100", 
"10000101", 
"10110101", 
"01101101", 
"10000100", 
"01000011", 
"01111111", 
"10000001", 
"10110110", 
"01110110", 
"01101111", 
"01111010", 
"10100100", 
"01110000", 
"10001111", 
"01010001", 
"10001101", 
"01111100", 
"01110100", 
"01111100", 
"10001110", 
"01100101", 
"01111001", 
"10010000", 
"01101100", 
"10111101", 
"01101110", 
"01101001", 
"10001100", 
"01111001", 
"10010110", 
"01110011", 
"01110100", 
"10010001", 
"10101100", 
"01111011", 
"10001001", 
"10000001", 
"01011000", 
"10001111", 
"10011000", 
"10100101", 
"10010000", 
"01101000", 
"10101010", 
"10100101", 
"01111110", 
"01111011", 
"10000100", 
"10000101", 
"01100001", 
"01111110", 
"01010110", 
"01110000", 
"01101100", 
"10000101", 
"10110110", 
"10010100", 
"10011010", 
"10010100", 
"10110110", 
"10001001", 
"10001101", 
"01010101", 
"01110010", 
"01111001", 
"10011000", 
"01110100", 
"10000111", 
"01100110", 
"01011111", 
"01101001", 
"10100100", 
"01011001", 
"01110010", 
"01100100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_84: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_84(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
