use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_101_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_101_LAYER;

architecture Behavioral of ROM_FC_120_101_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_101: ROM_ARRAY_PESOS_FC_120 := (
"10000110", 
"10011011", 
"01100000", 
"01100011", 
"10000000", 
"10001100", 
"01100000", 
"01101111", 
"10000111", 
"00111100", 
"01000100", 
"01110111", 
"01000010", 
"10101000", 
"01110010", 
"01110010", 
"10000010", 
"01100001", 
"01011001", 
"01100011", 
"10000001", 
"10110111", 
"01111101", 
"01011100", 
"10010110", 
"00111110", 
"10011101", 
"01001010", 
"01101100", 
"11000000", 
"01111011", 
"10001100", 
"10000100", 
"01100101", 
"01100000", 
"10011110", 
"01110001", 
"10001111", 
"10001010", 
"01101011", 
"01110111", 
"01110110", 
"10110101", 
"10000000", 
"01111010", 
"10101111", 
"10001010", 
"10001101", 
"01111111", 
"10000011", 
"10001011", 
"10001101", 
"01111111", 
"10000100", 
"10000101", 
"01110000", 
"10010110", 
"01111011", 
"10000010", 
"01111111", 
"01001111", 
"11000101", 
"10010001", 
"10001010", 
"10010000", 
"10101101", 
"01011100", 
"01111101", 
"01111111", 
"10000101", 
"01110011", 
"10000110", 
"10001110", 
"01011111", 
"01110111", 
"01101001", 
"01100111", 
"10000111", 
"10000010", 
"01110101", 
"10000010", 
"10000100", 
"01101101", 
"01000100", 
"01110011", 
"10100000", 
"10000111", 
"01110110", 
"01111001", 
"01101111", 
"10000010", 
"01100011", 
"01000110", 
"01100101", 
"10010010", 
"10000001", 
"01011010", 
"01100001", 
"01110100", 
"01101011", 
"01110010", 
"01110001", 
"10010011", 
"01011010", 
"10010001", 
"01101010", 
"10000100", 
"01101100", 
"01100000", 
"10010100", 
"01111100", 
"10001001", 
"01110010", 
"01011011", 
"01100111", 
"10100100", 
"10001101", 
"01110101", 
"01111000", 
"01010101", 
"10001000", 
"10010000", 
"01100110", 
"10001000", 
"01110001", 
"10010101", 
"01110100", 
"01110011", 
"10010010", 
"10001011", 
"01100000", 
"01011101", 
"10000100", 
"10010100", 
"01010101", 
"01010010", 
"10001100", 
"01011110", 
"10001010", 
"01101111", 
"01100110", 
"01110010", 
"01111100", 
"01110010", 
"10000110", 
"01100110", 
"01101000", 
"01100000", 
"10001100", 
"10110001", 
"01111011", 
"01011110", 
"10010010", 
"01101111", 
"10001100", 
"01010001", 
"01011100", 
"01010010", 
"10001011", 
"10001111", 
"10010011", 
"01100111", 
"10010101", 
"10001101", 
"10001101", 
"10011100", 
"10011111", 
"01011110", 
"10011101", 
"10000101", 
"01111001", 
"01101011", 
"01110110", 
"10011010", 
"10010011", 
"01111011", 
"01111001", 
"01010011", 
"01101100", 
"01100100", 
"01110001", 
"10000110", 
"10001001", 
"01101001", 
"10000110", 
"10010011", 
"01110111", 
"01110101", 
"10001101", 
"10001000", 
"10000111", 
"01110010", 
"10011010", 
"10000011", 
"01011110", 
"01110001", 
"10010011", 
"10100110", 
"01101101", 
"01100000", 
"10000111", 
"01111101", 
"10000000", 
"01111101", 
"01111110", 
"01010100", 
"10000011", 
"10010010", 
"01110011", 
"01101001", 
"01111101", 
"01100011", 
"10000110", 
"10010000", 
"01100000", 
"10000111", 
"10001010", 
"01100000", 
"01111101", 
"01111011", 
"01010001", 
"01101010", 
"10000011", 
"10000011", 
"10011100", 
"01110110", 
"01110010", 
"10001010", 
"01111011", 
"10001111", 
"10101001", 
"10010010", 
"10001000", 
"01100000", 
"10011000", 
"01110010", 
"01110011", 
"01111110", 
"01111011", 
"10000010", 
"10000110", 
"10000000", 
"01101000", 
"01111110", 
"01110000", 
"10010100", 
"10011011", 
"01101011", 
"01101011", 
"01001110", 
"10100001", 
"01110001", 
"10100101", 
"10001010", 
"10001011", 
"10010001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_101: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_101(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
