use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_40_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_40_LAYER;

architecture Behavioral of ROM_FC_84_40_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_40: ROM_ARRAY_PESOS_FC_84 := (
"01010100", 
"10001101", 
"01100111", 
"01101000", 
"01110011", 
"01110110", 
"10011011", 
"10000101", 
"01100100", 
"10010111", 
"10011000", 
"01101001", 
"01011111", 
"01010010", 
"01111100", 
"01100111", 
"10000011", 
"01111011", 
"01101100", 
"01110000", 
"10001010", 
"10100101", 
"10000011", 
"01110011", 
"01101000", 
"10010010", 
"01110011", 
"10000110", 
"01101010", 
"01011100", 
"01110010", 
"10001000", 
"01111101", 
"01101001", 
"10000111", 
"01010100", 
"10001101", 
"10000011", 
"01010110", 
"01101111", 
"10010000", 
"10101100", 
"01010111", 
"01110001", 
"01100101", 
"01111100", 
"01011110", 
"01111100", 
"01110101", 
"10001101", 
"01011010", 
"10000101", 
"01100101", 
"01101110", 
"01110101", 
"01110000", 
"01101010", 
"10011010", 
"01011100", 
"11001110", 
"10001100", 
"01100110", 
"01110100", 
"01100001", 
"10010011", 
"10011011", 
"01110111", 
"01101111", 
"01110001", 
"01110000", 
"10010101", 
"01100111", 
"01011000", 
"01111101", 
"10000100", 
"01110101", 
"10010111", 
"10001011", 
"01011111", 
"01011100", 
"10000011", 
"10000111", 
"01101111", 
"10010011", 
"01110010", 
"01101111", 
"10010110", 
"10000001", 
"01101101", 
"10010001", 
"01100110", 
"01110000", 
"10010100", 
"10000001", 
"01100010", 
"10010011", 
"01101001", 
"01111000", 
"01101000", 
"01100010", 
"10000110", 
"10000100", 
"01110100", 
"01111100", 
"01110001", 
"10000000", 
"10001011", 
"10000011", 
"01101100", 
"01110100", 
"01011100", 
"10011111", 
"01111010", 
"10001000", 
"10010110", 
"01101011", 
"10010000", 
"01101000", 
"01110110", 
"01101000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_40: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_40(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
