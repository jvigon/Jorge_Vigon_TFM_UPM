use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_110_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_110_LAYER;

architecture Behavioral of ROM_FC_120_110_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_110: ROM_ARRAY_PESOS_FC_120 := (
"01111110", 
"01010100", 
"10001100", 
"10010101", 
"01110110", 
"00110100", 
"10010000", 
"01100010", 
"01111010", 
"01110010", 
"01011101", 
"01101100", 
"10001001", 
"01001011", 
"01101111", 
"01110000", 
"01110011", 
"01101100", 
"10101111", 
"10010001", 
"01101100", 
"01011100", 
"10101000", 
"01111000", 
"01101100", 
"10001100", 
"10000000", 
"00101010", 
"01101011", 
"00110100", 
"10001100", 
"01110100", 
"01111111", 
"10101111", 
"10110000", 
"10110000", 
"01111000", 
"10000100", 
"01101010", 
"10001000", 
"01110000", 
"01010111", 
"10000100", 
"01111011", 
"01010100", 
"01101010", 
"10001000", 
"10001111", 
"10001011", 
"10110011", 
"01000101", 
"01100101", 
"01101001", 
"01011000", 
"01100011", 
"01100000", 
"10001110", 
"00010000", 
"01111100", 
"00100110", 
"01110110", 
"10010110", 
"10001000", 
"01100100", 
"01111010", 
"01000000", 
"10000000", 
"10101110", 
"01101100", 
"01010000", 
"01001010", 
"01011010", 
"01111011", 
"10010100", 
"01001111", 
"00000000", 
"00011110", 
"10101110", 
"01110000", 
"01110100", 
"01110110", 
"01011000", 
"01111110", 
"10000110", 
"01101101", 
"01111111", 
"01101010", 
"01111000", 
"01101011", 
"10110101", 
"01000101", 
"01010001", 
"10000110", 
"10000000", 
"01111011", 
"01111000", 
"01010111", 
"10111010", 
"10001001", 
"01111110", 
"01110000", 
"10111101", 
"01001100", 
"10001110", 
"10001100", 
"10101111", 
"01110110", 
"01110010", 
"10000110", 
"01111110", 
"01111110", 
"10001110", 
"01110110", 
"01101101", 
"10000110", 
"01010000", 
"10000100", 
"10101011", 
"10100110", 
"10100110", 
"01110100", 
"10000001", 
"10001111", 
"10010111", 
"01011000", 
"01100011", 
"01111110", 
"10000111", 
"10010100", 
"01100101", 
"01010110", 
"01100011", 
"01101100", 
"01011001", 
"01001000", 
"01111000", 
"10000011", 
"01111101", 
"01001111", 
"10001011", 
"01101011", 
"10001111", 
"01111011", 
"10000001", 
"01111111", 
"01111001", 
"01100110", 
"01101110", 
"01111111", 
"01010101", 
"01110111", 
"01111110", 
"10001110", 
"10101110", 
"01010101", 
"11010101", 
"10010000", 
"10011010", 
"10001010", 
"01110011", 
"01010010", 
"01011000", 
"01011101", 
"01001101", 
"10001110", 
"01101101", 
"01101010", 
"10010101", 
"01101110", 
"01100100", 
"01001000", 
"10001101", 
"01101111", 
"01100010", 
"10001101", 
"10000000", 
"10010001", 
"01110000", 
"10101001", 
"01110010", 
"10000101", 
"01011110", 
"10011100", 
"01111001", 
"01101101", 
"01111100", 
"01110101", 
"01000011", 
"01111011", 
"01100110", 
"10001010", 
"10000001", 
"10011010", 
"01111100", 
"10011110", 
"00100110", 
"01110011", 
"10001111", 
"01011010", 
"01101110", 
"01101101", 
"10010111", 
"10000011", 
"01000110", 
"10011001", 
"01111111", 
"10001000", 
"10000111", 
"10000101", 
"01010101", 
"10001111", 
"01101111", 
"01110101", 
"01101011", 
"10010001", 
"01111110", 
"01110111", 
"01011000", 
"10000010", 
"10000000", 
"10001011", 
"10101110", 
"10001111", 
"10000010", 
"10100100", 
"10010001", 
"10001000", 
"01010011", 
"10001000", 
"10000001", 
"01110001", 
"01100100", 
"01110000", 
"01111100", 
"01001100", 
"10000000", 
"10000100", 
"01110000", 
"01111001", 
"01110010", 
"10111101", 
"01011100", 
"10010010", 
"01010110", 
"10000011", 
"01101111", 
"11000100", 
"01100010", 
"10000011", 
"10001101", 
"01111001", 
"01000111", 
"01001000", 
"10001010", 
"01110010", 
"01111101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_110 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_110(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
