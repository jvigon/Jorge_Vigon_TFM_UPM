use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_69_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_69_LAYER;

architecture Behavioral of ROM_FC_84_69_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_69: ROM_ARRAY_PESOS_FC_84 := (
"01110100", 
"10000010", 
"01001010", 
"01111101", 
"01011110", 
"10000101", 
"01111010", 
"01110110", 
"01111110", 
"10001111", 
"10000101", 
"01001001", 
"01010001", 
"11100101", 
"10001110", 
"10000011", 
"01111000", 
"01101101", 
"01110101", 
"10001000", 
"01111101", 
"01011110", 
"01101001", 
"10000101", 
"10000010", 
"01110100", 
"01011110", 
"10000001", 
"10001100", 
"01011000", 
"01101101", 
"01010011", 
"10001101", 
"01111101", 
"01111111", 
"01011010", 
"01100001", 
"01110100", 
"01110101", 
"10010100", 
"10000111", 
"10001110", 
"01101011", 
"10000111", 
"01101001", 
"01100100", 
"10001011", 
"01110000", 
"01100011", 
"01111001", 
"01101001", 
"10011000", 
"10000111", 
"01100111", 
"01100000", 
"01100011", 
"10000011", 
"01110011", 
"10000110", 
"10000101", 
"01011011", 
"01111101", 
"10000010", 
"10001101", 
"01001011", 
"01100111", 
"10000110", 
"01110010", 
"10001110", 
"01111111", 
"01011000", 
"01101110", 
"01001111", 
"01011001", 
"10010000", 
"01110001", 
"10000110", 
"01110101", 
"10000100", 
"01100100", 
"10001011", 
"01101101", 
"01000011", 
"01010100", 
"01001011", 
"01101111", 
"01101101", 
"01111101", 
"01100101", 
"10000101", 
"01010010", 
"10000111", 
"01010010", 
"01111001", 
"01011100", 
"10000000", 
"01010101", 
"01101000", 
"01101001", 
"10000000", 
"01100111", 
"01001010", 
"01100101", 
"10000001", 
"01011010", 
"10000000", 
"01110010", 
"01110011", 
"01000011", 
"11000100", 
"01101010", 
"01111011", 
"01110111", 
"10000001", 
"10011001", 
"10001000", 
"01100000", 
"10101010", 
"01101010", 
"01001100"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_69: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_69(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
