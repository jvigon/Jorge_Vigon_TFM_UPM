use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_116_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_116_LAYER;

architecture Behavioral of ROM_FC_120_116_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_116: ROM_ARRAY_PESOS_FC_120 := (
"01111101", 
"01000111", 
"01111111", 
"10001000", 
"01111100", 
"00001101", 
"01110111", 
"10000111", 
"01110001", 
"10011010", 
"01011011", 
"01110011", 
"10010111", 
"01110101", 
"10010000", 
"01101110", 
"10010101", 
"01101001", 
"10000001", 
"10011110", 
"10101001", 
"01011000", 
"10100010", 
"01101010", 
"01110111", 
"10001111", 
"01001001", 
"10100111", 
"10100101", 
"00010110", 
"10010000", 
"01111011", 
"01111001", 
"01000001", 
"01111001", 
"10010001", 
"10011001", 
"10011001", 
"01011111", 
"10011101", 
"10010001", 
"10010001", 
"10001011", 
"10001110", 
"01101110", 
"01101011", 
"10001011", 
"01110100", 
"10010000", 
"10000001", 
"01110011", 
"10000001", 
"01111111", 
"10000011", 
"01110111", 
"10010111", 
"01111000", 
"01110011", 
"01111011", 
"01101011", 
"01011110", 
"01011100", 
"01110011", 
"10000110", 
"10000010", 
"10000100", 
"01011101", 
"01011001", 
"01110000", 
"01011100", 
"01110010", 
"01100000", 
"10001001", 
"10100010", 
"01111011", 
"01111100", 
"00011000", 
"10110011", 
"01111110", 
"10010001", 
"01010100", 
"01110000", 
"01110111", 
"10010001", 
"01111110", 
"01001110", 
"01111011", 
"01101000", 
"01111100", 
"10000100", 
"01100010", 
"01100001", 
"01011111", 
"01110110", 
"10011110", 
"10001001", 
"01011001", 
"01100010", 
"01110110", 
"01110100", 
"10000110", 
"10010111", 
"01000100", 
"01100100", 
"01111100", 
"01111101", 
"10000001", 
"01100010", 
"01111011", 
"10000010", 
"01110010", 
"10000110", 
"10000011", 
"01011111", 
"01101011", 
"01111011", 
"01111000", 
"01111110", 
"10101100", 
"10011101", 
"10001001", 
"10100100", 
"01011111", 
"01110010", 
"01101101", 
"01000011", 
"10010100", 
"01100011", 
"10100111", 
"01101001", 
"01111100", 
"10011000", 
"10001010", 
"01111010", 
"00010110", 
"01110110", 
"01111011", 
"01110110", 
"01110010", 
"10001110", 
"01101100", 
"10100000", 
"01111000", 
"01110100", 
"01110000", 
"01111100", 
"01101110", 
"10011010", 
"01011000", 
"01111011", 
"10000110", 
"01110110", 
"10000111", 
"10001010", 
"01011010", 
"01110001", 
"01101000", 
"10101100", 
"10011000", 
"01110110", 
"10000100", 
"01111000", 
"01001100", 
"10000001", 
"01110011", 
"11001010", 
"01001110", 
"10000110", 
"10100110", 
"10000100", 
"01110100", 
"01101001", 
"01101111", 
"01100001", 
"10010001", 
"01111011", 
"01110101", 
"01101001", 
"10100100", 
"10011001", 
"01111001", 
"01110101", 
"10011110", 
"01111100", 
"10011001", 
"01111011", 
"01111101", 
"01011010", 
"01000010", 
"10011010", 
"10010000", 
"10000100", 
"10011011", 
"01100110", 
"10100101", 
"01111010", 
"01111010", 
"01111101", 
"01110010", 
"01101111", 
"01111101", 
"01111100", 
"01001111", 
"01111110", 
"10001100", 
"01101110", 
"10011100", 
"10000111", 
"10000001", 
"01001000", 
"10010100", 
"01110000", 
"10001001", 
"01111000", 
"01110011", 
"01110101", 
"10001001", 
"10011101", 
"00111010", 
"01110010", 
"10100100", 
"01101000", 
"10001100", 
"10000011", 
"01010001", 
"01011001", 
"10001100", 
"10001011", 
"10000101", 
"10001101", 
"10000000", 
"01110011", 
"10001001", 
"10000100", 
"01111011", 
"10000001", 
"10010011", 
"10000101", 
"10010101", 
"10000101", 
"01100000", 
"01110001", 
"10011010", 
"10011101", 
"10000010", 
"01111110", 
"10011001", 
"01001111", 
"10000111", 
"01101111", 
"10001010", 
"01111000", 
"01000011", 
"01011010", 
"10010001", 
"10000011"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_116 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_116(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
