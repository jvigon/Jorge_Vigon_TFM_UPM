use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_70_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_70_LAYER;

architecture Behavioral of ROM_FC_120_70_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_70: ROM_ARRAY_PESOS_FC_120 := (
"10001001", 
"01110111", 
"10001110", 
"10101000", 
"01111101", 
"01111011", 
"01000111", 
"10000001", 
"01110111", 
"10010110", 
"01011100", 
"10001001", 
"01010100", 
"10111101", 
"10000000", 
"01110100", 
"10010010", 
"01000001", 
"01101110", 
"01111101", 
"10001110", 
"01111100", 
"01111101", 
"10001001", 
"10000011", 
"01110000", 
"01011000", 
"01111011", 
"01100000", 
"10101100", 
"10001101", 
"10101011", 
"10010001", 
"01111011", 
"10010100", 
"01110111", 
"01110011", 
"01101100", 
"10010100", 
"01110011", 
"01101111", 
"10001000", 
"10000001", 
"01011011", 
"01101000", 
"10101001", 
"10000100", 
"10010110", 
"01101100", 
"01100001", 
"10101000", 
"01110110", 
"10000110", 
"01010100", 
"10100001", 
"10100000", 
"10001011", 
"01100101", 
"01101000", 
"11001011", 
"10011011", 
"01101011", 
"10000011", 
"10011001", 
"01111101", 
"10111010", 
"01110011", 
"00011111", 
"01111000", 
"01111010", 
"10011010", 
"01111101", 
"10001011", 
"10000010", 
"10000000", 
"10001110", 
"10110100", 
"01000101", 
"10001110", 
"01111111", 
"01111010", 
"10011110", 
"01100110", 
"01010111", 
"01110010", 
"01111100", 
"01100001", 
"01110001", 
"01110010", 
"10001010", 
"01011001", 
"01110111", 
"01111101", 
"01110101", 
"10001011", 
"10000001", 
"01110011", 
"01110111", 
"01111111", 
"10001111", 
"10010011", 
"01101011", 
"01111111", 
"01101001", 
"10000000", 
"01101011", 
"01110101", 
"10000010", 
"10010011", 
"10000100", 
"10000111", 
"10000110", 
"01001011", 
"01100101", 
"10100011", 
"10000101", 
"10001110", 
"01010111", 
"01101101", 
"01100111", 
"10000000", 
"01100101", 
"01100011", 
"10000000", 
"10010111", 
"01010011", 
"10001001", 
"01110101", 
"10000110", 
"10000001", 
"10011010", 
"01101111", 
"01111110", 
"10100101", 
"10010111", 
"01110110", 
"10000011", 
"10001010", 
"10100010", 
"10010110", 
"10011000", 
"01100011", 
"01111110", 
"01110011", 
"01111010", 
"01111011", 
"01011101", 
"01011010", 
"01111100", 
"10011000", 
"01110001", 
"10100101", 
"01110110", 
"10000010", 
"01100110", 
"10000101", 
"01101000", 
"10000101", 
"10000000", 
"10000110", 
"01110000", 
"10100000", 
"01110001", 
"01010101", 
"01111011", 
"10001001", 
"10010001", 
"10000010", 
"01110110", 
"01100011", 
"01111110", 
"11010000", 
"10010010", 
"01101010", 
"10000110", 
"01110010", 
"01011011", 
"01110111", 
"01110101", 
"01000001", 
"01110011", 
"10001100", 
"10001010", 
"10001000", 
"10000110", 
"01111011", 
"01100001", 
"01101001", 
"01111011", 
"01011000", 
"10001010", 
"01110001", 
"01111011", 
"01101100", 
"01010101", 
"10101101", 
"01111101", 
"01111000", 
"10011001", 
"01110010", 
"10001001", 
"01100101", 
"10001011", 
"01100000", 
"00111111", 
"10001000", 
"10001010", 
"01111101", 
"01101110", 
"01011110", 
"01110110", 
"10001111", 
"10000000", 
"10001010", 
"10010011", 
"01111000", 
"10000111", 
"01010001", 
"01110111", 
"01111001", 
"01010101", 
"10100101", 
"10001001", 
"01110000", 
"01110011", 
"01001010", 
"01111111", 
"01011111", 
"10001111", 
"10000100", 
"10100101", 
"01111001", 
"10000011", 
"01100110", 
"01101101", 
"10010111", 
"10000100", 
"01101101", 
"01110110", 
"01111011", 
"10000011", 
"10000010", 
"01100111", 
"01110001", 
"10010000", 
"10000010", 
"10010100", 
"10010110", 
"01110010", 
"01011011", 
"01111000", 
"01101110", 
"01101001", 
"01010101", 
"10000101", 
"10001000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_70: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_70(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
