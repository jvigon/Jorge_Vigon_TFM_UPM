use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_119_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_119_LAYER;

architecture Behavioral of ROM_FC_120_119_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_119: ROM_ARRAY_PESOS_FC_120 := (
"10101010", 
"01101100", 
"01101101", 
"00100111", 
"10101000", 
"01010001", 
"00101110", 
"01100011", 
"01111010", 
"10010101", 
"10000001", 
"10101110", 
"10010101", 
"01111000", 
"10001011", 
"10010111", 
"01100010", 
"01110111", 
"01110100", 
"01000101", 
"10011011", 
"10010000", 
"01001011", 
"01101101", 
"10010010", 
"01110100", 
"01111100", 
"10010011", 
"01100000", 
"10001101", 
"10000110", 
"10001111", 
"10100100", 
"10101101", 
"01111011", 
"01010010", 
"10010010", 
"10100111", 
"01101010", 
"01110011", 
"01110110", 
"01101001", 
"01110010", 
"10101001", 
"01011001", 
"11010100", 
"10100101", 
"10010010", 
"10010100", 
"10010011", 
"01000000", 
"10001101", 
"01100110", 
"10000000", 
"01100001", 
"10010001", 
"10001010", 
"00100111", 
"01110110", 
"01110000", 
"01011101", 
"11000001", 
"10101001", 
"10000010", 
"10100000", 
"01111110", 
"10100111", 
"00110111", 
"01100001", 
"01000100", 
"01111011", 
"11011001", 
"10010011", 
"10011101", 
"00111111", 
"10011000", 
"10011010", 
"10110011", 
"10000110", 
"10011100", 
"01110011", 
"10000011", 
"01110110", 
"01001100", 
"01101001", 
"10010001", 
"01011101", 
"11000011", 
"01111011", 
"01011010", 
"01100000", 
"10100010", 
"10011110", 
"10010000", 
"10000000", 
"10010011", 
"10100001", 
"01101101", 
"01011001", 
"01101001", 
"10000000", 
"01111001", 
"01111101", 
"10010110", 
"10000000", 
"01110101", 
"01101100", 
"10010110", 
"10110010", 
"11000000", 
"10010011", 
"10000000", 
"10010010", 
"01111000", 
"10101111", 
"10000100", 
"01110100", 
"10010110", 
"10011001", 
"10000111", 
"01110100", 
"01100100", 
"01011110", 
"10001001", 
"10001010", 
"01111110", 
"10000100", 
"01110100", 
"01011100", 
"01100111", 
"10011000", 
"01001011", 
"10101110", 
"01111000", 
"11000010", 
"10100011", 
"01101011", 
"10000000", 
"01110001", 
"01111110", 
"10111011", 
"10011101", 
"10000101", 
"10011101", 
"10100011", 
"10001100", 
"10011101", 
"01100001", 
"10010010", 
"10000111", 
"10011011", 
"01111100", 
"10001011", 
"10011101", 
"01011010", 
"10010010", 
"10010001", 
"01011000", 
"01111111", 
"10001010", 
"01111101", 
"10010010", 
"01111000", 
"10001101", 
"01111011", 
"00110001", 
"01101011", 
"10000101", 
"10010010", 
"01110011", 
"10000111", 
"01101000", 
"10000000", 
"10001101", 
"01110111", 
"10011100", 
"10000010", 
"01101100", 
"10000010", 
"10010011", 
"01111010", 
"01000110", 
"01100111", 
"01110000", 
"10010111", 
"10100110", 
"10011010", 
"01110110", 
"10011011", 
"01101101", 
"10010110", 
"10001001", 
"01110101", 
"01011010", 
"10001110", 
"01110001", 
"01111001", 
"01110111", 
"01111100", 
"10011000", 
"01111000", 
"01111100", 
"10110000", 
"01001001", 
"10000100", 
"01110010", 
"01111000", 
"10001000", 
"01011010", 
"10100010", 
"10101111", 
"01111011", 
"10000100", 
"01100010", 
"01101010", 
"10100011", 
"01101110", 
"10011001", 
"01111000", 
"01110001", 
"10111000", 
"01010110", 
"10000001", 
"10010111", 
"10001111", 
"10110110", 
"10011001", 
"10000101", 
"10000100", 
"01101010", 
"01110001", 
"10001110", 
"10001110", 
"10001100", 
"01011001", 
"10101000", 
"01101110", 
"01111100", 
"10000010", 
"10000011", 
"00110011", 
"01011011", 
"10001111", 
"11001110", 
"10001000", 
"01110001", 
"00100111", 
"01100010", 
"01111001", 
"10110011", 
"01100101", 
"11000100", 
"10011110", 
"10010001", 
"10001110", 
"10000010"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_119 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_119(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
