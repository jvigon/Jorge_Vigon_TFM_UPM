use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_115_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_115_LAYER;

architecture Behavioral of ROM_FC_120_115_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_115: ROM_ARRAY_PESOS_FC_120 := (
"01110000", 
"10000111", 
"01011100", 
"01101001", 
"01111111", 
"01000001", 
"01110110", 
"10000000", 
"01111100", 
"10100101", 
"01110001", 
"10111100", 
"01100110", 
"01110011", 
"10000000", 
"10001011", 
"01001001", 
"10000000", 
"01100100", 
"00111101", 
"10001111", 
"01100110", 
"01101010", 
"01111011", 
"10000101", 
"10001011", 
"10111010", 
"10011101", 
"10010000", 
"00111100", 
"10100111", 
"10100001", 
"01100011", 
"01110111", 
"01011010", 
"00100001", 
"10001011", 
"01111111", 
"01110000", 
"01110100", 
"10000111", 
"01000101", 
"10011100", 
"10001000", 
"01001001", 
"10101100", 
"10100010", 
"10101010", 
"01100101", 
"01011100", 
"01011001", 
"01101000", 
"10010000", 
"01111010", 
"01111110", 
"01111110", 
"10010001", 
"10000001", 
"01101101", 
"01110011", 
"10100000", 
"11010010", 
"10011000", 
"10001101", 
"10100000", 
"01111000", 
"01010101", 
"01101101", 
"01011011", 
"10011100", 
"01111010", 
"10001101", 
"01100100", 
"01101000", 
"01011010", 
"01111000", 
"10001000", 
"01010010", 
"10001101", 
"10001100", 
"10011101", 
"01011111", 
"01101101", 
"01011011", 
"01110010", 
"10010000", 
"01100100", 
"01011001", 
"01101100", 
"01011100", 
"01100110", 
"10010110", 
"01111010", 
"11001010", 
"10001110", 
"10000001", 
"10001110", 
"10001110", 
"01100110", 
"01101110", 
"10001100", 
"01110100", 
"10000010", 
"01111100", 
"10000010", 
"01001011", 
"01111111", 
"01100100", 
"01001110", 
"10100010", 
"10001010", 
"01110111", 
"01110111", 
"01010100", 
"01010010", 
"01101101", 
"01111010", 
"01111111", 
"01101110", 
"01010100", 
"10010101", 
"01100111", 
"10001010", 
"10100000", 
"10000100", 
"10010000", 
"01101101", 
"10000010", 
"01100010", 
"01111101", 
"01010100", 
"01100000", 
"10001111", 
"10000011", 
"01111100", 
"10010111", 
"10000111", 
"01011110", 
"01011100", 
"00101011", 
"10000100", 
"01110010", 
"10000001", 
"01110100", 
"10100011", 
"01111011", 
"01101110", 
"01110111", 
"10001001", 
"10000111", 
"10001010", 
"10010011", 
"10001110", 
"01011010", 
"01101110", 
"01101001", 
"01110111", 
"10011101", 
"01111101", 
"01111110", 
"10001010", 
"01101101", 
"01111010", 
"01001000", 
"10001101", 
"01100101", 
"01110011", 
"01110100", 
"10100110", 
"01011001", 
"01001100", 
"01010000", 
"01111111", 
"10010011", 
"01111011", 
"01111111", 
"10011111", 
"01101110", 
"01101111", 
"00111101", 
"01111110", 
"10000100", 
"01101111", 
"01110101", 
"10100110", 
"01110111", 
"01110110", 
"10000010", 
"10001111", 
"00100110", 
"10001100", 
"01111010", 
"01110000", 
"01111000", 
"10000100", 
"10000001", 
"01100010", 
"01100111", 
"10001010", 
"01110110", 
"10001101", 
"01101000", 
"10010001", 
"01011001", 
"01100010", 
"01101100", 
"10010010", 
"10001101", 
"01100101", 
"10011010", 
"10001100", 
"10001001", 
"10010010", 
"01111101", 
"10000001", 
"01100000", 
"10011001", 
"01011000", 
"01110110", 
"01100100", 
"01100110", 
"01101100", 
"01111001", 
"10011011", 
"01101100", 
"10000010", 
"10110010", 
"10100010", 
"01110100", 
"01100111", 
"01011111", 
"01100111", 
"10100100", 
"10000100", 
"10000010", 
"01110100", 
"10000110", 
"01011010", 
"01110110", 
"01111001", 
"01110100", 
"10001001", 
"10101001", 
"01110011", 
"10001100", 
"01111000", 
"01000101", 
"10010110", 
"10011111", 
"01111111", 
"01111011", 
"10000110", 
"10100000", 
"01011011", 
"10010111", 
"01110110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_115 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_115(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
