use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_46_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_46_LAYER;

architecture Behavioral of ROM_FC_120_46_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_46: ROM_ARRAY_PESOS_FC_120 := (
"01110011", 
"01100001", 
"01010000", 
"10001101", 
"01011010", 
"01001011", 
"01101110", 
"01011010", 
"01101111", 
"00110110", 
"10000011", 
"01100010", 
"10000111", 
"01101000", 
"10000001", 
"10000010", 
"00011110", 
"01111001", 
"01101110", 
"01000110", 
"10011011", 
"01111100", 
"01110100", 
"01010110", 
"01111101", 
"01011011", 
"10100111", 
"10010101", 
"10011010", 
"01101010", 
"10010101", 
"01100010", 
"00010110", 
"10001110", 
"10011110", 
"01111100", 
"01110000", 
"00110000", 
"01010100", 
"01100111", 
"01111010", 
"10111110", 
"01100000", 
"01010010", 
"10010010", 
"01000101", 
"01110001", 
"10000001", 
"00111100", 
"10000000", 
"01110011", 
"01100101", 
"01101001", 
"01111010", 
"01111101", 
"01010010", 
"01111000", 
"10001000", 
"01110011", 
"11000000", 
"10011010", 
"10000010", 
"01111100", 
"10000111", 
"01100000", 
"10111110", 
"01101001", 
"01101011", 
"10000100", 
"10010110", 
"01111011", 
"01011111", 
"01101000", 
"00101101", 
"10000100", 
"01111101", 
"10010011", 
"00000110", 
"10000110", 
"10000101", 
"01110011", 
"10001001", 
"01110110", 
"01110000", 
"01011010", 
"10001010", 
"10101110", 
"01001111", 
"01110001", 
"00100111", 
"01101000", 
"01001100", 
"10011101", 
"01100110", 
"10010101", 
"01110101", 
"01110000", 
"10010011", 
"10011111", 
"01110011", 
"01101110", 
"01010111", 
"01110010", 
"10010010", 
"10000111", 
"01010001", 
"01101011", 
"01010001", 
"10010100", 
"11100111", 
"01110111", 
"10000101", 
"10001101", 
"10011011", 
"10001001", 
"01000110", 
"10000010", 
"01111101", 
"10011101", 
"01111101", 
"01101011", 
"10110110", 
"01100011", 
"10011010", 
"10000101", 
"01101001", 
"01100011", 
"10010100", 
"10010101", 
"10010101", 
"10001011", 
"01111001", 
"10100001", 
"10111011", 
"10101100", 
"01110111", 
"01110101", 
"00101101", 
"10000111", 
"10101111", 
"10010111", 
"00110001", 
"10000111", 
"01101010", 
"01101100", 
"10101010", 
"01001000", 
"01110110", 
"01010101", 
"10001011", 
"10000001", 
"01110100", 
"01111011", 
"01011111", 
"10000000", 
"01001111", 
"01110000", 
"01100111", 
"01110100", 
"10000100", 
"01100001", 
"01100011", 
"10000111", 
"01101011", 
"01101001", 
"10010110", 
"10110111", 
"01101010", 
"01110101", 
"01101111", 
"10110000", 
"10100011", 
"10000101", 
"10000111", 
"01110011", 
"01100001", 
"10001101", 
"01110101", 
"00100011", 
"01100011", 
"01101101", 
"10000000", 
"10010101", 
"10000110", 
"10001111", 
"01111111", 
"01001111", 
"01110001", 
"01000111", 
"01101111", 
"10000011", 
"01101110", 
"01100111", 
"01010001", 
"10011001", 
"10011101", 
"10110011", 
"01101011", 
"01010001", 
"01000100", 
"01111100", 
"10001100", 
"01101111", 
"00111110", 
"10011011", 
"00011000", 
"10000110", 
"01111010", 
"00111111", 
"01011111", 
"10101011", 
"10100110", 
"01101111", 
"01011001", 
"10011101", 
"01101110", 
"10011100", 
"10010110", 
"10001101", 
"01000111", 
"01111101", 
"10100010", 
"01111100", 
"01111100", 
"01111111", 
"00111010", 
"10110101", 
"01110000", 
"01101111", 
"10000010", 
"01111111", 
"10001010", 
"01110101", 
"10010110", 
"01100111", 
"10000111", 
"10000100", 
"01010100", 
"01111010", 
"10011010", 
"10011100", 
"01111010", 
"00011101", 
"00010011", 
"10010101", 
"01111101", 
"10110111", 
"10111000", 
"10010011", 
"01110001", 
"01010001", 
"01000110", 
"01101111", 
"10000001", 
"10001000", 
"01110111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_46: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_46(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
