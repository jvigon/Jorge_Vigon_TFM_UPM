use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_80_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_80_LAYER;

architecture Behavioral of ROM_FC_84_80_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_80: ROM_ARRAY_PESOS_FC_84 := (
"01111010", 
"10000000", 
"01100001", 
"01110100", 
"10010101", 
"01111110", 
"10010110", 
"10001111", 
"10100011", 
"01110110", 
"01100100", 
"01100000", 
"10001111", 
"01110010", 
"00110001", 
"01100111", 
"01110010", 
"01111000", 
"01101110", 
"10001010", 
"01110110", 
"10110101", 
"10010101", 
"01111100", 
"10010011", 
"01110111", 
"10000011", 
"01110100", 
"10000010", 
"01100101", 
"10010111", 
"10001010", 
"01101001", 
"10100001", 
"01111101", 
"01000110", 
"10011111", 
"01111100", 
"01111010", 
"01010010", 
"10001001", 
"10010010", 
"10100000", 
"10001011", 
"00101110", 
"01111011", 
"01010001", 
"10010001", 
"10001100", 
"10000111", 
"01000110", 
"10000011", 
"10010110", 
"01101000", 
"10011110", 
"10100000", 
"01101011", 
"01100110", 
"10000010", 
"10101000", 
"10010010", 
"01110100", 
"01011001", 
"10011111", 
"01110001", 
"01110101", 
"10100110", 
"10000001", 
"01111010", 
"10001101", 
"01101100", 
"01111100", 
"01000111", 
"10110001", 
"10000000", 
"01100110", 
"10110001", 
"01110111", 
"01011010", 
"01111000", 
"10111101", 
"01111011", 
"01110000", 
"01101111", 
"01111101", 
"01111100", 
"10000011", 
"10011000", 
"10010011", 
"10000111", 
"01100100", 
"10100111", 
"01111000", 
"10001011", 
"10001110", 
"01110100", 
"01101110", 
"01111001", 
"01001000", 
"01010000", 
"01111111", 
"01101111", 
"01110000", 
"10011001", 
"10011100", 
"01111110", 
"01111010", 
"01110110", 
"01111111", 
"10101111", 
"10010010", 
"10000101", 
"10000001", 
"10000101", 
"10001101", 
"10001111", 
"01000111", 
"10000001", 
"10001010", 
"10010101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_80: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_80(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
