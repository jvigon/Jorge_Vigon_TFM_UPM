use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_89_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_89_LAYER;

architecture Behavioral of ROM_FC_120_89_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_89: ROM_ARRAY_PESOS_FC_120 := (
"10001011", 
"10100101", 
"10000010", 
"01000000", 
"01011101", 
"01001111", 
"10100010", 
"01111101", 
"01111001", 
"01101001", 
"01010111", 
"00111001", 
"10010100", 
"01011110", 
"01111100", 
"10000111", 
"01010011", 
"10001001", 
"01110100", 
"00010010", 
"01110111", 
"01001001", 
"10111001", 
"10000010", 
"01111101", 
"10010000", 
"10000101", 
"01111100", 
"10011010", 
"01000100", 
"10001000", 
"01111110", 
"00111111", 
"10000010", 
"01010111", 
"01001000", 
"10000110", 
"01110111", 
"01101111", 
"10000001", 
"01110001", 
"10000001", 
"10100011", 
"10000001", 
"10001011", 
"10001111", 
"10010001", 
"01111010", 
"01010001", 
"01111011", 
"01100011", 
"01111010", 
"01111000", 
"10011111", 
"10000011", 
"01011010", 
"01110110", 
"00101001", 
"10001100", 
"01101000", 
"01110101", 
"10011000", 
"01110100", 
"10001100", 
"10001100", 
"10100010", 
"01101001", 
"10001011", 
"01100100", 
"10101110", 
"10001111", 
"01101010", 
"10000011", 
"01011000", 
"10011011", 
"01101101", 
"01110101", 
"01001111", 
"10001111", 
"01111010", 
"01110011", 
"10010110", 
"10011110", 
"00101111", 
"10000010", 
"10001111", 
"01100001", 
"00110010", 
"01111000", 
"10000000", 
"10100011", 
"01100111", 
"00111100", 
"01000101", 
"10010010", 
"01110110", 
"01111000", 
"10010100", 
"10100111", 
"01010110", 
"10000011", 
"10000011", 
"01111000", 
"01011100", 
"10000110", 
"01001000", 
"10001011", 
"10000001", 
"01010000", 
"10011100", 
"10000011", 
"10010100", 
"01101110", 
"10101111", 
"01011110", 
"01111001", 
"10010101", 
"10000111", 
"10101000", 
"01010100", 
"10000011", 
"01011110", 
"10000010", 
"01111001", 
"01100010", 
"01111101", 
"01111111", 
"01101111", 
"10001101", 
"10000100", 
"01011110", 
"10000000", 
"10010001", 
"10101001", 
"01101010", 
"10101000", 
"10100011", 
"01100000", 
"10101111", 
"01011001", 
"00011111", 
"10110100", 
"01101010", 
"01101111", 
"01111100", 
"01011101", 
"01110101", 
"01101110", 
"10001100", 
"10010100", 
"10110110", 
"01111111", 
"10101101", 
"01001111", 
"10010000", 
"10000010", 
"00011001", 
"10101100", 
"01111111", 
"01101111", 
"01101111", 
"01011001", 
"10001000", 
"10011100", 
"01111110", 
"10000111", 
"10010101", 
"10001111", 
"10001000", 
"00110011", 
"01100110", 
"10100000", 
"01010011", 
"10010001", 
"01111100", 
"01100101", 
"10101001", 
"01010001", 
"01000011", 
"00010001", 
"10001100", 
"01110101", 
"10011111", 
"01101001", 
"01111110", 
"01101010", 
"01110100", 
"10001111", 
"01111101", 
"01001010", 
"10010001", 
"10000001", 
"10100011", 
"01010111", 
"10100010", 
"10011111", 
"01110010", 
"10110001", 
"10000011", 
"10010111", 
"01111100", 
"00110001", 
"10001001", 
"00000000", 
"01011010", 
"01110011", 
"01110101", 
"10001111", 
"01101111", 
"00101011", 
"10110101", 
"10111000", 
"01101110", 
"10001111", 
"10011000", 
"01001111", 
"10001100", 
"01100100", 
"01100011", 
"01011010", 
"01100000", 
"10110110", 
"10010000", 
"01110111", 
"10001001", 
"01100011", 
"10111011", 
"10011101", 
"01111001", 
"10010000", 
"10010110", 
"10001010", 
"01111000", 
"10011001", 
"01101011", 
"01010010", 
"10100101", 
"10000000", 
"01110000", 
"01111101", 
"10011110", 
"01100011", 
"10010010", 
"10000001", 
"10010010", 
"01100101", 
"10000101", 
"10011111", 
"01101000", 
"10000100", 
"01101110", 
"01000011", 
"01111110", 
"01001100", 
"10001100", 
"01111110"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_89: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_89(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
