use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_43_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_43_LAYER;

architecture Behavioral of ROM_FC_84_43_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_43: ROM_ARRAY_PESOS_FC_84 := (
"01110001", 
"10001110", 
"10001111", 
"10000100", 
"01101100", 
"01101111", 
"10001100", 
"10001110", 
"01111100", 
"01111000", 
"01110101", 
"01100000", 
"01011000", 
"01010100", 
"11001011", 
"01011000", 
"01000000", 
"01011110", 
"01101001", 
"10001000", 
"01101110", 
"01101010", 
"10100011", 
"01110111", 
"01111010", 
"10010111", 
"01000000", 
"01101111", 
"01010011", 
"01101111", 
"10001101", 
"10001110", 
"01110101", 
"10010110", 
"10000010", 
"01010111", 
"10110000", 
"01110011", 
"01100011", 
"01111001", 
"01111011", 
"01110010", 
"10001001", 
"01101101", 
"01011101", 
"01111111", 
"01101001", 
"10010000", 
"01100000", 
"01101111", 
"01110110", 
"10000001", 
"10001101", 
"01111000", 
"01011011", 
"10010001", 
"10001010", 
"10000110", 
"10010010", 
"10001011", 
"01101111", 
"01100110", 
"01101011", 
"01111100", 
"01101110", 
"01111011", 
"01111000", 
"10010010", 
"10001000", 
"10000111", 
"10100011", 
"01100110", 
"01000000", 
"01000101", 
"01100110", 
"01111101", 
"10010110", 
"01001111", 
"01100011", 
"10001111", 
"01011110", 
"10000001", 
"01011110", 
"01011011", 
"01011111", 
"01010111", 
"01111011", 
"01000011", 
"01101111", 
"01100110", 
"01100111", 
"10001111", 
"01101110", 
"01111110", 
"01110000", 
"10001011", 
"01010110", 
"10010101", 
"01101110", 
"01110100", 
"10010010", 
"01100001", 
"01100011", 
"00110011", 
"01100010", 
"01101000", 
"10001001", 
"10000101", 
"01111011", 
"11001001", 
"01000101", 
"01101001", 
"01110001", 
"01111110", 
"10010000", 
"01011001", 
"01100100", 
"00111101", 
"10000010", 
"01111001"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_43: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_43(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
