use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_58_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_58_LAYER;

architecture Behavioral of ROM_FC_120_58_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_58: ROM_ARRAY_PESOS_FC_120 := (
"01111011", 
"01111010", 
"10000001", 
"10100011", 
"01101110", 
"10001101", 
"10001110", 
"01010001", 
"10001100", 
"01000111", 
"10010110", 
"00101000", 
"01011101", 
"10110010", 
"10000000", 
"10000100", 
"01111000", 
"01011000", 
"10000001", 
"10010110", 
"01110000", 
"01110000", 
"10001010", 
"01110111", 
"01110111", 
"10010111", 
"10011000", 
"01000001", 
"01101101", 
"10000010", 
"01101010", 
"10001100", 
"01111000", 
"01100010", 
"01101110", 
"10000010", 
"01111100", 
"00111101", 
"00111110", 
"01101100", 
"10001000", 
"10011100", 
"01110001", 
"01100101", 
"01101100", 
"01010111", 
"10000100", 
"10000100", 
"01011000", 
"01000101", 
"10000011", 
"01101101", 
"01110000", 
"01111010", 
"01010101", 
"10010001", 
"01110110", 
"10100101", 
"01011001", 
"10010110", 
"10000000", 
"01101110", 
"10000000", 
"01100000", 
"01100011", 
"10100011", 
"01111011", 
"01000111", 
"01100100", 
"10011001", 
"01110100", 
"01010101", 
"01101111", 
"10011110", 
"10011011", 
"01000110", 
"01111010", 
"00101111", 
"10000011", 
"01111110", 
"10000011", 
"10011000", 
"01110110", 
"01101010", 
"01110000", 
"01111100", 
"01100011", 
"01010110", 
"10001111", 
"10011101", 
"10011101", 
"10000100", 
"01101110", 
"01111011", 
"01110111", 
"10000011", 
"01100110", 
"10000100", 
"01111011", 
"01101000", 
"10010001", 
"01100111", 
"01100100", 
"01001110", 
"10000110", 
"10001111", 
"01110110", 
"10000111", 
"10011000", 
"10001100", 
"10000111", 
"10001010", 
"01110101", 
"10011010", 
"01100000", 
"00011111", 
"10001010", 
"01111011", 
"01110110", 
"01000110", 
"10001010", 
"10000110", 
"10000010", 
"10011100", 
"10100111", 
"01110100", 
"01111000", 
"10000001", 
"10000001", 
"01110000", 
"10010101", 
"01100111", 
"01111110", 
"10011111", 
"01010111", 
"10111010", 
"01110110", 
"10100010", 
"01111111", 
"10000001", 
"10000101", 
"10001110", 
"10001011", 
"10010000", 
"10000011", 
"01110000", 
"01100010", 
"00111111", 
"01110011", 
"10010110", 
"01111010", 
"10000111", 
"01101011", 
"10011111", 
"01101111", 
"10011000", 
"01100111", 
"01111111", 
"01110010", 
"01111011", 
"10100100", 
"10100110", 
"01010111", 
"01001111", 
"01110101", 
"10001101", 
"01111011", 
"10000000", 
"10000001", 
"01110000", 
"01100000", 
"10101110", 
"01101011", 
"10011110", 
"10000101", 
"10000001", 
"10011101", 
"10001111", 
"10000101", 
"00011101", 
"01110000", 
"10001010", 
"10110001", 
"01101101", 
"10010010", 
"01001011", 
"10000100", 
"11000100", 
"10100010", 
"01111101", 
"10010100", 
"10010100", 
"10000101", 
"01110011", 
"01100110", 
"01100110", 
"01110101", 
"01101100", 
"01110111", 
"10100101", 
"10001010", 
"01110100", 
"10010010", 
"01110100", 
"10000010", 
"10010000", 
"01110100", 
"01111101", 
"10010010", 
"10000011", 
"10001000", 
"10000101", 
"10010010", 
"01110010", 
"01101001", 
"10010010", 
"01101110", 
"01010011", 
"01011011", 
"10000110", 
"10001010", 
"01111000", 
"10001111", 
"10010100", 
"10011010", 
"10101011", 
"01111001", 
"01010011", 
"10010000", 
"10010011", 
"10101110", 
"01111000", 
"01101101", 
"01010011", 
"01110010", 
"10010011", 
"10000001", 
"10010110", 
"01111011", 
"10000110", 
"10010001", 
"10001010", 
"01111010", 
"01000111", 
"10001110", 
"10000011", 
"01110000", 
"01100110", 
"10010100", 
"01100011", 
"10001001", 
"10001100", 
"10101010", 
"10001110", 
"10001000", 
"10000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_58: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_58(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
