use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_67_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_67_LAYER;

architecture Behavioral of ROM_FC_84_67_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_67: ROM_ARRAY_PESOS_FC_84 := (
"01100100", 
"01100010", 
"01111110", 
"10001110", 
"10000001", 
"10010010", 
"01111101", 
"10001010", 
"01101001", 
"01101001", 
"01111010", 
"01110110", 
"01110110", 
"01110110", 
"10001101", 
"01011111", 
"01100111", 
"01110010", 
"01100001", 
"10000101", 
"01011110", 
"01111000", 
"10001111", 
"01110110", 
"01111111", 
"01110101", 
"10001111", 
"01101010", 
"01100100", 
"01100111", 
"10000011", 
"01101100", 
"10011000", 
"10010011", 
"10001010", 
"01010101", 
"10001000", 
"01110011", 
"10000111", 
"01111101", 
"01110110", 
"01111001", 
"01111000", 
"01100001", 
"01100001", 
"10000010", 
"01100110", 
"10010100", 
"10001010", 
"10000000", 
"10001110", 
"01101110", 
"10001101", 
"01101011", 
"10000010", 
"10001110", 
"10000100", 
"10001001", 
"01101100", 
"10001001", 
"10001001", 
"01110010", 
"10001000", 
"01110011", 
"01100101", 
"10001111", 
"01111001", 
"01101110", 
"01110000", 
"10011011", 
"10000110", 
"01101001", 
"10001000", 
"01100110", 
"01110101", 
"10010001", 
"10011100", 
"10000110", 
"01100000", 
"01101000", 
"10000100", 
"01011111", 
"10000001", 
"01100011", 
"01010011", 
"01101010", 
"01110101", 
"01010101", 
"10000000", 
"01101010", 
"01110111", 
"10000100", 
"10001101", 
"10000101", 
"01101001", 
"01111100", 
"01111111", 
"01101001", 
"10001000", 
"01110110", 
"10010111", 
"10001111", 
"10000110", 
"01100110", 
"01101111", 
"01101010", 
"10000110", 
"10010010", 
"01100111", 
"01111101", 
"10001010", 
"10000101", 
"01101111", 
"01110111", 
"01110110", 
"10000011", 
"10000100", 
"01101011", 
"10000011", 
"01100101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_67: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_67(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
