use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_56_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_56_LAYER;

architecture Behavioral of ROM_FC_84_56_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_84_56: ROM_ARRAY_PESOS_FC_84 := (
"01001101", 
"10010101", 
"10011011", 
"01100111", 
"00111001", 
"01011111", 
"10011001", 
"01110101", 
"01011111", 
"01010111", 
"01111101", 
"00110111", 
"01011110", 
"01101111", 
"10000110", 
"10000001", 
"01000101", 
"10110101", 
"00111111", 
"00101100", 
"10010101", 
"01110110", 
"01100100", 
"10001101", 
"01100101", 
"10011000", 
"10001001", 
"10001001", 
"10000111", 
"10000101", 
"01110111", 
"10011000", 
"10100101", 
"10100000", 
"10000001", 
"10100011", 
"10001010", 
"01001101", 
"01000101", 
"01111110", 
"00100011", 
"11011011", 
"01111100", 
"00111000", 
"01011000", 
"01011000", 
"10001011", 
"10100000", 
"01111000", 
"01101011", 
"01100100", 
"10011000", 
"10010110", 
"10011100", 
"01111001", 
"10101010", 
"10000010", 
"01101110", 
"01011011", 
"11001011", 
"01110001", 
"01101101", 
"10101001", 
"01010101", 
"01110100", 
"01110011", 
"01101010", 
"10111110", 
"10010110", 
"01011001", 
"10010101", 
"00101101", 
"01111001", 
"10000010", 
"01110111", 
"01110100", 
"01101001", 
"01100101", 
"10100001", 
"01001100", 
"01001111", 
"01111010", 
"01111110", 
"10010100", 
"01010011", 
"10000000", 
"01000011", 
"10010001", 
"10011000", 
"01111110", 
"01101011", 
"10010110", 
"10001000", 
"01011000", 
"10010100", 
"10000101", 
"10010001", 
"10010000", 
"01111010", 
"01001111", 
"01110111", 
"10110110", 
"01000000", 
"01011101", 
"10000000", 
"01110010", 
"10001001", 
"01011011", 
"01111011", 
"11000101", 
"01100000", 
"10010000", 
"01100101", 
"10001110", 
"01110111", 
"01100110", 
"10010001", 
"10001010", 
"10000100", 
"01011000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_56 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_56(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
