use work.Package_FC_84.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_84_51_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC_84)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_84_51_LAYER;

architecture Behavioral of ROM_FC_84_51_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_84 is Array (0 to (Dim_pesos_FC_84-1)) of STD_LOGIC_VECTOR(7 downto 0);
signal ROM_FC_84_51: ROM_ARRAY_PESOS_FC_84 := (
"01110101", 
"01100010", 
"10000100", 
"01100100", 
"10111100", 
"10010101", 
"01101101", 
"10011101", 
"10010101", 
"01011011", 
"10011110", 
"10100000", 
"01101010", 
"10000011", 
"10100011", 
"01110101", 
"10001101", 
"10010010", 
"10011110", 
"01111000", 
"10111010", 
"10011011", 
"10010110", 
"01101101", 
"10000101", 
"10010110", 
"10001000", 
"10010011", 
"10100101", 
"01011011", 
"10010101", 
"01110010", 
"01101100", 
"01111010", 
"00101110", 
"01101001", 
"01101000", 
"01110000", 
"10011001", 
"01011011", 
"10101001", 
"10001100", 
"10000111", 
"01100111", 
"10000010", 
"01011011", 
"01010111", 
"01011011", 
"10010011", 
"01111011", 
"10000111", 
"10001101", 
"10010000", 
"01100100", 
"10011110", 
"01110001", 
"10000111", 
"01110001", 
"10100001", 
"01010100", 
"10100001", 
"10000010", 
"01111001", 
"10100011", 
"01001110", 
"10000011", 
"10000001", 
"10010101", 
"01110000", 
"01100110", 
"01111101", 
"10110110", 
"01110000", 
"01111000", 
"01111001", 
"10000100", 
"10001011", 
"01100011", 
"10000001", 
"10000101", 
"01110111", 
"10100110", 
"01101000", 
"01011001", 
"10011011", 
"10000100", 
"01110100", 
"10001001", 
"01101000", 
"01110010", 
"10010001", 
"01101110", 
"10000010", 
"01011010", 
"01111010", 
"10000100", 
"01101000", 
"10000101", 
"10100001", 
"10000010", 
"01110000", 
"01111110", 
"01100101", 
"01101110", 
"10011010", 
"10010001", 
"01110001", 
"10000110", 
"01001000", 
"01010011", 
"10011100", 
"01110101", 
"01110001", 
"01111000", 
"10001100", 
"10000011", 
"10000011", 
"01110001", 
"10000110", 
"01011111"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_84_51: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_84_51(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
