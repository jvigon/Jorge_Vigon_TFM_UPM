use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_50_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_50_LAYER;

architecture Behavioral of ROM_FC_120_50_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_50: ROM_ARRAY_PESOS_FC_120 := (
"10100111", 
"10100001", 
"11000000", 
"10010011", 
"10000000", 
"10101101", 
"01111000", 
"01111000", 
"01111110", 
"01111010", 
"01101000", 
"00110111", 
"01101100", 
"11000110", 
"01101101", 
"10011011", 
"10010111", 
"01111110", 
"01000110", 
"01001011", 
"01011010", 
"10010000", 
"10001100", 
"10000010", 
"10010110", 
"01111100", 
"01110011", 
"00110001", 
"10010000", 
"10100100", 
"01111010", 
"01110111", 
"10000100", 
"01100101", 
"01111011", 
"10000001", 
"10010000", 
"01100000", 
"01101011", 
"01010111", 
"01101110", 
"01110111", 
"01101001", 
"01000011", 
"01111110", 
"10110001", 
"01100110", 
"10000101", 
"01100110", 
"01100000", 
"10111010", 
"01101001", 
"01111110", 
"10110011", 
"01101010", 
"01110101", 
"10000111", 
"01111010", 
"01000100", 
"01010011", 
"01111000", 
"01111101", 
"01111111", 
"10001101", 
"01111000", 
"01111111", 
"01010101", 
"01101001", 
"10000011", 
"10101010", 
"01111011", 
"01111100", 
"10001101", 
"10110110", 
"10100110", 
"01111001", 
"10101001", 
"01001011", 
"10000101", 
"01101001", 
"10011000", 
"10011011", 
"01100110", 
"00111001", 
"01111010", 
"10010010", 
"01110001", 
"10001110", 
"01111011", 
"10010011", 
"10101100", 
"10110001", 
"01110001", 
"00111111", 
"01111010", 
"10000111", 
"01110110", 
"10001011", 
"10010000", 
"01110000", 
"01111110", 
"01000010", 
"10000111", 
"01011000", 
"01110011", 
"10100001", 
"01111000", 
"10011001", 
"01011100", 
"01110011", 
"10000101", 
"10001010", 
"01110000", 
"10111011", 
"01010111", 
"01100011", 
"01110110", 
"10000100", 
"00101111", 
"10010010", 
"10001111", 
"10011100", 
"10010010", 
"10011110", 
"01101111", 
"01111010", 
"10000011", 
"10000110", 
"01110111", 
"01110010", 
"10000001", 
"01010011", 
"10010111", 
"01111001", 
"01100100", 
"11001100", 
"01110100", 
"10000100", 
"10001011", 
"01001011", 
"01100001", 
"10000111", 
"01111101", 
"01111110", 
"01111001", 
"01101010", 
"01101011", 
"01010010", 
"10000011", 
"10000010", 
"10000110", 
"10011010", 
"01100111", 
"01000010", 
"01111010", 
"10010001", 
"01011000", 
"10101010", 
"01010110", 
"01110110", 
"10100100", 
"01011101", 
"01110111", 
"01111000", 
"10001011", 
"10011000", 
"10100010", 
"01110011", 
"10001110", 
"01100101", 
"01010011", 
"10000001", 
"00111011", 
"10001000", 
"01111101", 
"10000100", 
"10101101", 
"10010011", 
"01101111", 
"01110011", 
"01111101", 
"10101010", 
"01111100", 
"10010100", 
"10011010", 
"00111001", 
"01101111", 
"10100011", 
"10010110", 
"10000110", 
"01110011", 
"01111101", 
"01100001", 
"01100000", 
"01011111", 
"01000110", 
"10000001", 
"01111011", 
"10011010", 
"10111011", 
"10000101", 
"01100000", 
"01011110", 
"01001010", 
"00111011", 
"10001001", 
"01101111", 
"10010011", 
"10001101", 
"01100001", 
"01010010", 
"01100000", 
"01110101", 
"01111100", 
"10011010", 
"01110110", 
"01111111", 
"01010101", 
"01011001", 
"01000110", 
"01001001", 
"00111100", 
"10000101", 
"01111011", 
"10100011", 
"01001100", 
"01010001", 
"01111110", 
"10001111", 
"10010010", 
"10010101", 
"01111001", 
"10001101", 
"01110111", 
"01110000", 
"01100110", 
"01100000", 
"01101111", 
"10000011", 
"01111100", 
"01110010", 
"01001111", 
"01000101", 
"10100000", 
"01110010", 
"01101010", 
"01001001", 
"10000100", 
"10100010", 
"01100011", 
"10011000", 
"01011111", 
"01100011", 
"01100110", 
"10001000", 
"10001101"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_50: signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_50(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
