use work.Package_FC_120.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity ROM_FC_120_108_LAYER is
        Port ( CLK : in STD_LOGIC;
           addra_pool_2 : IN STD_LOGIC_VECTOR((log2c(Dim_pesos_FC)-1) downto 0);
           douta_pool_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
           );
end ROM_FC_120_108_LAYER;

architecture Behavioral of ROM_FC_120_108_LAYER is
--SIGNAL W_next, W_reg : STD_LOGIC_VECTOR(7 DOWNTO 0);
TYPE ROM_ARRAY_PESOS_FC_120 is Array (0 to (Dim_pesos_FC-1)) of STD_LOGIC_VECTOR(7 downto 0);--2400 16 filtros de 5x5x6
signal ROM_FC_120_108: ROM_ARRAY_PESOS_FC_120 := (
"01101011", 
"01110111", 
"10011101", 
"01011011", 
"10001101", 
"01001010", 
"01011011", 
"01100111", 
"01111000", 
"10101101", 
"01111011", 
"10001001", 
"10001110", 
"10010111", 
"10000111", 
"10001101", 
"10001100", 
"10010010", 
"01110001", 
"01110101", 
"10111110", 
"01010010", 
"10000101", 
"01110001", 
"01101110", 
"10100001", 
"01111101", 
"01101100", 
"10000111", 
"01010111", 
"10000000", 
"10010000", 
"01111000", 
"10011000", 
"01111010", 
"01111101", 
"10000011", 
"10000000", 
"01110111", 
"01010010", 
"10000010", 
"01110100", 
"01111110", 
"10010010", 
"10000010", 
"01111011", 
"10000110", 
"01110111", 
"01111110", 
"10000001", 
"10010101", 
"01100110", 
"10010111", 
"10011011", 
"10000100", 
"01011011", 
"10100101", 
"01001001", 
"01111110", 
"10101011", 
"10110011", 
"10010110", 
"10010100", 
"01110101", 
"10100000", 
"10010101", 
"01111111", 
"01100010", 
"11001001", 
"01111011", 
"10010001", 
"10110000", 
"01011001", 
"10100000", 
"10010100", 
"01111101", 
"01100001", 
"10010110", 
"01110111", 
"01101101", 
"10010111", 
"10000001", 
"01010011", 
"01000100", 
"10001011", 
"01111000", 
"01001110", 
"01111000", 
"01110101", 
"10000111", 
"01001101", 
"10001001", 
"01100010", 
"10100100", 
"01111010", 
"10000010", 
"10110001", 
"10001011", 
"01000101", 
"00100011", 
"01011100", 
"01111100", 
"10010110", 
"10001000", 
"01011100", 
"01111110", 
"01111010", 
"10011010", 
"01110011", 
"10000010", 
"10001011", 
"01101110", 
"10010100", 
"10000111", 
"01100010", 
"00111101", 
"01100100", 
"10011110", 
"10111001", 
"01101101", 
"10100101", 
"01110100", 
"10010101", 
"11001000", 
"01101111", 
"10000101", 
"01100001", 
"10001001", 
"10011101", 
"01100111", 
"10001001", 
"01001111", 
"10110010", 
"10001001", 
"10111110", 
"10111000", 
"01110101", 
"01011000", 
"10010101", 
"01111111", 
"10010011", 
"01111101", 
"01111001", 
"01101011", 
"11001011", 
"10010010", 
"01010111", 
"01111001", 
"01100001", 
"10010100", 
"01111101", 
"10101101", 
"10000111", 
"01010110", 
"01011100", 
"10010011", 
"10011001", 
"10100011", 
"10001110", 
"10001100", 
"10011101", 
"01000101", 
"01111100", 
"01111110", 
"01100101", 
"01000000", 
"10100101", 
"11000000", 
"01110101", 
"01000001", 
"00110101", 
"01100111", 
"10000001", 
"01001111", 
"01110111", 
"01110000", 
"10011010", 
"01000000", 
"01111101", 
"01110110", 
"10001001", 
"01101011", 
"10010010", 
"01111010", 
"10101001", 
"10001010", 
"01101000", 
"01001001", 
"01110111", 
"01101000", 
"01111100", 
"01101011", 
"01100011", 
"01001001", 
"10010110", 
"10010011", 
"01100010", 
"10010100", 
"10001110", 
"01110011", 
"01110001", 
"10010001", 
"10111000", 
"01010111", 
"10010010", 
"00010010", 
"10000110", 
"01111111", 
"01100011", 
"10001111", 
"01110000", 
"10001011", 
"01100000", 
"01101000", 
"01010001", 
"10010110", 
"01110010", 
"10010110", 
"10011011", 
"10001000", 
"10011011", 
"01111101", 
"10001001", 
"10010001", 
"01001000", 
"01100011", 
"10110111", 
"10100100", 
"01111111", 
"00110101", 
"10000000", 
"01111000", 
"10011101", 
"10101010", 
"01011001", 
"01011110", 
"01111000", 
"01000100", 
"10001100", 
"10000101", 
"01000100", 
"00010100", 
"10100011", 
"10111000", 
"10000111", 
"00111100", 
"00000000", 
"01101111", 
"10010110", 
"10111100", 
"01001001", 
"10010110", 
"10011001", 
"01011100", 
"01111011", 
"10000000"
);
attribute rom_style : string;
attribute rom_style of ROM_FC_120_108 : signal is "block";
begin
   -- W_next <= ROM_FC_120_0(to_integer(unsigned(addra_pool_2)));
    --douta_pool_2 <= W_reg;

--    PROCESS (clk, reset)
--    BEGIN
--        IF reset = '0' THEN
--            W_reg <= (others => '0');
--        ELSIF CLK'event and CLK = '1' THEN
--            W_reg <= W_next;
--        END IF;
--    end process;

process(clk)
begin
if rising_edge(clk) then
    douta_pool_2<= ROM_FC_120_108(conv_integer(addra_pool_2));
end if;
end process;
end Behavioral;
